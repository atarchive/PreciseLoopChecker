// Gate Level Verilog Code Generated!
// GateLvl:500 GateNum:500 GateInputNum:2
// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_300, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_328, w_000_330, w_000_331, w_000_332, w_000_335, w_000_336, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_356, w_000_358, w_000_359, w_000_360, w_000_363, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_420, w_000_422, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_431, w_000_433, w_000_434, w_000_437, w_000_439, w_000_440, w_000_444, w_000_445, w_000_447, w_000_448, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_457, w_000_458, w_000_462, w_000_463, w_000_468, w_000_474, w_000_490, w_500_000, w_500_001, w_500_002, w_500_003, w_500_004, w_500_005, w_500_006, w_500_007, w_500_008, w_500_009, w_500_010, w_500_011, w_500_012, w_500_013, w_500_014, w_500_015, w_500_016, w_500_017, w_500_018, w_500_019, w_500_020, w_500_021, w_500_022, w_500_023, w_500_024, w_500_025, w_500_026, w_500_027, w_500_028, w_500_029, w_500_030, w_500_031, w_500_032, w_500_033, w_500_034, w_500_035, w_500_036, w_500_037, w_500_038, w_500_039, w_500_040, w_500_041, w_500_042, w_500_043, w_500_044, w_500_045, w_500_046, w_500_047, w_500_048, w_500_049, w_500_050, w_500_051, w_500_052, w_500_053, w_500_054, w_500_055, w_500_056, w_500_057, w_500_058, w_500_059, w_500_060, w_500_061, w_500_062, w_500_063, w_500_064, w_500_065, w_500_066, w_500_067, w_500_068, w_500_069, w_500_070, w_500_071, w_500_072, w_500_073, w_500_074, w_500_075, w_500_076, w_500_077, w_500_078, w_500_079, w_500_080, w_500_081, w_500_082, w_500_083, w_500_084, w_500_085, w_500_086, w_500_087, w_500_088, w_500_089, w_500_090, w_500_091, w_500_092, w_500_093, w_500_094, w_500_095, w_500_096, w_500_097, w_500_098, w_500_099, w_500_100, w_500_101, w_500_102, w_500_103, w_500_104, w_500_105, w_500_106, w_500_107, w_500_108, w_500_109, w_500_110, w_500_111, w_500_112, w_500_113, w_500_114, w_500_115, w_500_116, w_500_117, w_500_118, w_500_119, w_500_120, w_500_121, w_500_122, w_500_123, w_500_124, w_500_125, w_500_126, w_500_127, w_500_128, w_500_129, w_500_130, w_500_131, w_500_132, w_500_133, w_500_134, w_500_135, w_500_136, w_500_137, w_500_138, w_500_139, w_500_140, w_500_141, w_500_142, w_500_143, w_500_144, w_500_145, w_500_146, w_500_147, w_500_148, w_500_149, w_500_150, w_500_151, w_500_152, w_500_153, w_500_154, w_500_155, w_500_156, w_500_157, w_500_158, w_500_159, w_500_160, w_500_161, w_500_162, w_500_163, w_500_164, w_500_165, w_500_166, w_500_167, w_500_168, w_500_169, w_500_170, w_500_171, w_500_172, w_500_173, w_500_174, w_500_175, w_500_176, w_500_177, w_500_178, w_500_179, w_500_180, w_500_181, w_500_182, w_500_183, w_500_184, w_500_185, w_500_186, w_500_187, w_500_188, w_500_189, w_500_190, w_500_191, w_500_192, w_500_193, w_500_194, w_500_195, w_500_196, w_500_197, w_500_198, w_500_199, w_500_200, w_500_201, w_500_202, w_500_203, w_500_204, w_500_205, w_500_206, w_500_207, w_500_208, w_500_209, w_500_210, w_500_211, w_500_212, w_500_213, w_500_214, w_500_215, w_500_216, w_500_217, w_500_218, w_500_219, w_500_220, w_500_221, w_500_222, w_500_223, w_500_224, w_500_225, w_500_226, w_500_227, w_500_228, w_500_229, w_500_230, w_500_231, w_500_232, w_500_233, w_500_234, w_500_235, w_500_236, w_500_237, w_500_238, w_500_239, w_500_240, w_500_241, w_500_242, w_500_243, w_500_244, w_500_245, w_500_246, w_500_247, w_500_248, w_500_249, w_500_250, w_500_251, w_500_252, w_500_253, w_500_254, w_500_255, w_500_256, w_500_257, w_500_258, w_500_259, w_500_260, w_500_261, w_500_262, w_500_263, w_500_264, w_500_265, w_500_266, w_500_267, w_500_268, w_500_269, w_500_270, w_500_271, w_500_272, w_500_273, w_500_274, w_500_275, w_500_276, w_500_277, w_500_278, w_500_279, w_500_280, w_500_281, w_500_282, w_500_283, w_500_284, w_500_285, w_500_286, w_500_287, w_500_288, w_500_289, w_500_290, w_500_291, w_500_292, w_500_293, w_500_294, w_500_295, w_500_296, w_500_297, w_500_298, w_500_299, w_500_300, w_500_301, w_500_302, w_500_303, w_500_304, w_500_305, w_500_306, w_500_307, w_500_308, w_500_309, w_500_310, w_500_311, w_500_312, w_500_313, w_500_314, w_500_315, w_500_316, w_500_317, w_500_318, w_500_319, w_500_320, w_500_321, w_500_322, w_500_323, w_500_324, w_500_325, w_500_326, w_500_327, w_500_328, w_500_329, w_500_330, w_500_331, w_500_332, w_500_333, w_500_334, w_500_335, w_500_336, w_500_337, w_500_338, w_500_339, w_500_340, w_500_341, w_500_342, w_500_343, w_500_344, w_500_345, w_500_346, w_500_347, w_500_348, w_500_349, w_500_350, w_500_351, w_500_352, w_500_353, w_500_354, w_500_355, w_500_356, w_500_357, w_500_358, w_500_359, w_500_360, w_500_361, w_500_362, w_500_363, w_500_364, w_500_365, w_500_366, w_500_367, w_500_368, w_500_369, w_500_370, w_500_371, w_500_372, w_500_373, w_500_374, w_500_375, w_500_376, w_500_377, w_500_378, w_500_379, w_500_380, w_500_381, w_500_382, w_500_383, w_500_384, w_500_385, w_500_386, w_500_387, w_500_388, w_500_389, w_500_390, w_500_391, w_500_392, w_500_393, w_500_394, w_500_395, w_500_396, w_500_397, w_500_398, w_500_399, w_500_400, w_500_401, w_500_402, w_500_403, w_500_404, w_500_405, w_500_406, w_500_407, w_500_408, w_500_409, w_500_410, w_500_411, w_500_412, w_500_413, w_500_414, w_500_415, w_500_416, w_500_417, w_500_418, w_500_419, w_500_420, w_500_421, w_500_422, w_500_423, w_500_424, w_500_425, w_500_426, w_500_427, w_500_428, w_500_429, w_500_430, w_500_431, w_500_432, w_500_433, w_500_434, w_500_435, w_500_436, w_500_437, w_500_438, w_500_439, w_500_440, w_500_441, w_500_442, w_500_443, w_500_444, w_500_445, w_500_446, w_500_447, w_500_448, w_500_449, w_500_450, w_500_451, w_500_452, w_500_453, w_500_454, w_500_455, w_500_456, w_500_457, w_500_458, w_500_459, w_500_460, w_500_461, w_500_462, w_500_463, w_500_464 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_300, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_328, w_000_330, w_000_331, w_000_332, w_000_335, w_000_336, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_356, w_000_358, w_000_359, w_000_360, w_000_363, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_420, w_000_422, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_431, w_000_433, w_000_434, w_000_437, w_000_439, w_000_440, w_000_444, w_000_445, w_000_447, w_000_448, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_457, w_000_458, w_000_462, w_000_463, w_000_468, w_000_474, w_000_490;
  output w_500_000, w_500_001, w_500_002, w_500_003, w_500_004, w_500_005, w_500_006, w_500_007, w_500_008, w_500_009, w_500_010, w_500_011, w_500_012, w_500_013, w_500_014, w_500_015, w_500_016, w_500_017, w_500_018, w_500_019, w_500_020, w_500_021, w_500_022, w_500_023, w_500_024, w_500_025, w_500_026, w_500_027, w_500_028, w_500_029, w_500_030, w_500_031, w_500_032, w_500_033, w_500_034, w_500_035, w_500_036, w_500_037, w_500_038, w_500_039, w_500_040, w_500_041, w_500_042, w_500_043, w_500_044, w_500_045, w_500_046, w_500_047, w_500_048, w_500_049, w_500_050, w_500_051, w_500_052, w_500_053, w_500_054, w_500_055, w_500_056, w_500_057, w_500_058, w_500_059, w_500_060, w_500_061, w_500_062, w_500_063, w_500_064, w_500_065, w_500_066, w_500_067, w_500_068, w_500_069, w_500_070, w_500_071, w_500_072, w_500_073, w_500_074, w_500_075, w_500_076, w_500_077, w_500_078, w_500_079, w_500_080, w_500_081, w_500_082, w_500_083, w_500_084, w_500_085, w_500_086, w_500_087, w_500_088, w_500_089, w_500_090, w_500_091, w_500_092, w_500_093, w_500_094, w_500_095, w_500_096, w_500_097, w_500_098, w_500_099, w_500_100, w_500_101, w_500_102, w_500_103, w_500_104, w_500_105, w_500_106, w_500_107, w_500_108, w_500_109, w_500_110, w_500_111, w_500_112, w_500_113, w_500_114, w_500_115, w_500_116, w_500_117, w_500_118, w_500_119, w_500_120, w_500_121, w_500_122, w_500_123, w_500_124, w_500_125, w_500_126, w_500_127, w_500_128, w_500_129, w_500_130, w_500_131, w_500_132, w_500_133, w_500_134, w_500_135, w_500_136, w_500_137, w_500_138, w_500_139, w_500_140, w_500_141, w_500_142, w_500_143, w_500_144, w_500_145, w_500_146, w_500_147, w_500_148, w_500_149, w_500_150, w_500_151, w_500_152, w_500_153, w_500_154, w_500_155, w_500_156, w_500_157, w_500_158, w_500_159, w_500_160, w_500_161, w_500_162, w_500_163, w_500_164, w_500_165, w_500_166, w_500_167, w_500_168, w_500_169, w_500_170, w_500_171, w_500_172, w_500_173, w_500_174, w_500_175, w_500_176, w_500_177, w_500_178, w_500_179, w_500_180, w_500_181, w_500_182, w_500_183, w_500_184, w_500_185, w_500_186, w_500_187, w_500_188, w_500_189, w_500_190, w_500_191, w_500_192, w_500_193, w_500_194, w_500_195, w_500_196, w_500_197, w_500_198, w_500_199, w_500_200, w_500_201, w_500_202, w_500_203, w_500_204, w_500_205, w_500_206, w_500_207, w_500_208, w_500_209, w_500_210, w_500_211, w_500_212, w_500_213, w_500_214, w_500_215, w_500_216, w_500_217, w_500_218, w_500_219, w_500_220, w_500_221, w_500_222, w_500_223, w_500_224, w_500_225, w_500_226, w_500_227, w_500_228, w_500_229, w_500_230, w_500_231, w_500_232, w_500_233, w_500_234, w_500_235, w_500_236, w_500_237, w_500_238, w_500_239, w_500_240, w_500_241, w_500_242, w_500_243, w_500_244, w_500_245, w_500_246, w_500_247, w_500_248, w_500_249, w_500_250, w_500_251, w_500_252, w_500_253, w_500_254, w_500_255, w_500_256, w_500_257, w_500_258, w_500_259, w_500_260, w_500_261, w_500_262, w_500_263, w_500_264, w_500_265, w_500_266, w_500_267, w_500_268, w_500_269, w_500_270, w_500_271, w_500_272, w_500_273, w_500_274, w_500_275, w_500_276, w_500_277, w_500_278, w_500_279, w_500_280, w_500_281, w_500_282, w_500_283, w_500_284, w_500_285, w_500_286, w_500_287, w_500_288, w_500_289, w_500_290, w_500_291, w_500_292, w_500_293, w_500_294, w_500_295, w_500_296, w_500_297, w_500_298, w_500_299, w_500_300, w_500_301, w_500_302, w_500_303, w_500_304, w_500_305, w_500_306, w_500_307, w_500_308, w_500_309, w_500_310, w_500_311, w_500_312, w_500_313, w_500_314, w_500_315, w_500_316, w_500_317, w_500_318, w_500_319, w_500_320, w_500_321, w_500_322, w_500_323, w_500_324, w_500_325, w_500_326, w_500_327, w_500_328, w_500_329, w_500_330, w_500_331, w_500_332, w_500_333, w_500_334, w_500_335, w_500_336, w_500_337, w_500_338, w_500_339, w_500_340, w_500_341, w_500_342, w_500_343, w_500_344, w_500_345, w_500_346, w_500_347, w_500_348, w_500_349, w_500_350, w_500_351, w_500_352, w_500_353, w_500_354, w_500_355, w_500_356, w_500_357, w_500_358, w_500_359, w_500_360, w_500_361, w_500_362, w_500_363, w_500_364, w_500_365, w_500_366, w_500_367, w_500_368, w_500_369, w_500_370, w_500_371, w_500_372, w_500_373, w_500_374, w_500_375, w_500_376, w_500_377, w_500_378, w_500_379, w_500_380, w_500_381, w_500_382, w_500_383, w_500_384, w_500_385, w_500_386, w_500_387, w_500_388, w_500_389, w_500_390, w_500_391, w_500_392, w_500_393, w_500_394, w_500_395, w_500_396, w_500_397, w_500_398, w_500_399, w_500_400, w_500_401, w_500_402, w_500_403, w_500_404, w_500_405, w_500_406, w_500_407, w_500_408, w_500_409, w_500_410, w_500_411, w_500_412, w_500_413, w_500_414, w_500_415, w_500_416, w_500_417, w_500_418, w_500_419, w_500_420, w_500_421, w_500_422, w_500_423, w_500_424, w_500_425, w_500_426, w_500_427, w_500_428, w_500_429, w_500_430, w_500_431, w_500_432, w_500_433, w_500_434, w_500_435, w_500_436, w_500_437, w_500_438, w_500_439, w_500_440, w_500_441, w_500_442, w_500_443, w_500_444, w_500_445, w_500_446, w_500_447, w_500_448, w_500_449, w_500_450, w_500_451, w_500_452, w_500_453, w_500_454, w_500_455, w_500_456, w_500_457, w_500_458, w_500_459, w_500_460, w_500_461, w_500_462, w_500_463, w_500_464;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_300, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_328, w_000_330, w_000_331, w_000_332, w_000_335, w_000_336, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_356, w_000_358, w_000_359, w_000_360, w_000_363, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_420, w_000_422, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_431, w_000_433, w_000_434, w_000_437, w_000_439, w_000_440, w_000_444, w_000_445, w_000_447, w_000_448, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_457, w_000_458, w_000_462, w_000_463, w_000_468, w_000_474, w_000_490;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007, w_002_008, w_002_009, w_002_010, w_002_011, w_002_012, w_002_013, w_002_014, w_002_015, w_002_016, w_002_017, w_002_018, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_024, w_002_025, w_002_026, w_002_027;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023, w_003_024, w_003_025, w_003_026, w_003_027, w_003_028, w_003_029, w_003_030, w_003_031, w_003_032, w_003_033, w_003_034, w_003_035, w_003_036, w_003_037, w_003_038, w_003_039, w_003_040, w_003_041, w_003_042, w_003_043, w_003_044, w_003_045, w_003_046, w_003_047, w_003_048, w_003_049, w_003_050, w_003_051, w_003_052, w_003_053, w_003_054, w_003_055, w_003_056, w_003_057, w_003_058, w_003_059, w_003_060, w_003_061, w_003_062, w_003_063, w_003_064, w_003_065, w_003_066, w_003_067, w_003_068, w_003_069, w_003_070, w_003_071, w_003_072, w_003_073, w_003_074, w_003_075, w_003_076, w_003_077, w_003_078, w_003_079, w_003_080, w_003_081, w_003_082, w_003_083, w_003_084, w_003_085, w_003_086, w_003_087, w_003_088, w_003_089, w_003_090, w_003_091, w_003_092, w_003_093, w_003_094, w_003_095, w_003_096, w_003_097, w_003_098, w_003_099, w_003_100, w_003_101;
  wire w_004_000, w_004_001, w_004_002, w_004_003, w_004_004, w_004_005, w_004_006, w_004_007, w_004_008, w_004_009, w_004_010, w_004_011, w_004_012, w_004_014, w_004_015, w_004_016, w_004_017, w_004_018, w_004_019, w_004_020, w_004_021, w_004_022, w_004_023, w_004_024, w_004_025, w_004_026, w_004_027, w_004_028, w_004_029, w_004_030, w_004_031, w_004_032, w_004_034, w_004_036, w_004_037, w_004_038, w_004_039, w_004_043, w_004_044, w_004_046, w_004_047, w_004_048, w_004_050, w_004_051, w_004_052, w_004_053, w_004_054, w_004_057, w_004_058, w_004_059, w_004_060, w_004_061, w_004_062, w_004_065, w_004_066, w_004_067, w_004_069, w_004_070, w_004_071, w_004_072, w_004_076, w_004_078, w_004_080, w_004_081, w_004_082, w_004_083, w_004_084, w_004_085, w_004_086, w_004_087, w_004_088, w_004_089, w_004_091, w_004_094, w_004_095, w_004_096, w_004_097, w_004_098, w_004_100, w_004_102, w_004_103, w_004_104, w_004_105, w_004_106, w_004_107, w_004_109, w_004_110, w_004_111, w_004_112, w_004_113, w_004_114, w_004_115, w_004_117, w_004_118, w_004_120, w_004_121, w_004_122, w_004_124, w_004_125, w_004_127, w_004_128, w_004_130, w_004_131, w_004_132, w_004_133, w_004_134, w_004_135, w_004_136, w_004_137, w_004_138, w_004_139, w_004_141, w_004_142, w_004_143, w_004_144, w_004_147, w_004_148, w_004_149, w_004_152, w_004_154, w_004_155, w_004_156, w_004_157, w_004_159, w_004_160, w_004_161, w_004_163, w_004_164, w_004_166, w_004_167, w_004_168, w_004_172, w_004_173, w_004_175, w_004_178, w_004_179, w_004_180, w_004_181, w_004_182, w_004_183, w_004_184, w_004_186, w_004_187, w_004_188, w_004_189, w_004_190, w_004_191, w_004_192, w_004_193, w_004_194, w_004_195, w_004_198, w_004_199, w_004_201, w_004_202, w_004_203, w_004_204, w_004_206, w_004_209, w_004_210, w_004_211, w_004_213, w_004_214, w_004_215, w_004_216, w_004_217, w_004_219, w_004_221, w_004_222, w_004_223, w_004_224, w_004_225, w_004_226, w_004_227, w_004_228, w_004_230, w_004_232, w_004_233, w_004_234, w_004_237, w_004_238, w_004_239, w_004_240, w_004_241, w_004_243, w_004_244, w_004_245, w_004_246, w_004_247, w_004_249, w_004_250, w_004_251, w_004_252, w_004_253, w_004_254, w_004_255, w_004_256, w_004_257, w_004_259, w_004_260, w_004_263, w_004_265, w_004_267, w_004_268, w_004_269, w_004_271, w_004_272, w_004_273, w_004_274, w_004_275, w_004_276, w_004_277, w_004_278, w_004_279, w_004_280, w_004_282, w_004_283, w_004_285, w_004_286, w_004_287, w_004_289, w_004_290, w_004_291, w_004_292, w_004_293, w_004_295, w_004_296, w_004_297, w_004_300, w_004_301, w_004_302, w_004_303, w_004_304, w_004_305, w_004_307, w_004_308, w_004_309, w_004_310, w_004_311, w_004_312, w_004_313, w_004_314, w_004_315, w_004_316, w_004_317, w_004_318, w_004_319, w_004_320, w_004_321, w_004_322, w_004_323, w_004_324, w_004_325, w_004_327, w_004_328, w_004_329, w_004_330, w_004_331, w_004_332, w_004_333, w_004_336, w_004_338, w_004_339, w_004_340, w_004_341, w_004_342, w_004_343, w_004_344, w_004_345, w_004_346, w_004_347, w_004_348, w_004_349, w_004_350, w_004_351, w_004_352, w_004_353, w_004_354, w_004_356, w_004_357, w_004_358, w_004_359, w_004_360, w_004_361, w_004_362, w_004_363, w_004_365, w_004_366, w_004_367, w_004_368, w_004_369, w_004_370, w_004_371, w_004_372, w_004_373, w_004_374, w_004_376, w_004_378, w_004_380, w_004_381, w_004_383, w_004_384, w_004_385, w_004_386, w_004_387, w_004_388, w_004_389, w_004_393, w_004_394, w_004_395, w_004_396, w_004_397, w_004_398, w_004_399, w_004_400, w_004_401, w_004_402, w_004_405, w_004_406, w_004_407, w_004_408, w_004_410, w_004_412, w_004_413, w_004_415, w_004_416, w_004_417, w_004_418, w_004_419, w_004_421, w_004_424, w_004_425, w_004_426, w_004_427, w_004_428, w_004_429, w_004_430, w_004_431, w_004_432, w_004_433, w_004_435, w_004_436, w_004_438, w_004_439, w_004_440, w_004_441, w_004_442, w_004_444, w_004_445, w_004_446, w_004_447, w_004_448, w_004_449, w_004_451, w_004_452, w_004_454, w_004_455, w_004_456, w_004_457, w_004_458, w_004_459, w_004_460, w_004_462, w_004_463, w_004_464, w_004_465, w_004_467, w_004_468, w_004_469, w_004_470, w_004_471, w_004_472, w_004_473, w_004_474;
  wire w_005_000, w_005_001, w_005_002, w_005_003, w_005_004, w_005_005, w_005_006, w_005_007, w_005_008, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_017, w_005_018, w_005_019, w_005_020, w_005_021, w_005_022, w_005_023, w_005_024, w_005_025, w_005_026, w_005_027, w_005_028, w_005_029, w_005_030, w_005_031, w_005_032, w_005_033, w_005_034, w_005_035, w_005_036, w_005_037, w_005_038, w_005_039, w_005_040, w_005_041, w_005_042, w_005_043, w_005_044, w_005_045, w_005_046, w_005_047, w_005_048, w_005_049, w_005_050, w_005_052, w_005_053, w_005_055, w_005_056, w_005_057, w_005_058, w_005_059, w_005_060, w_005_061, w_005_062, w_005_064, w_005_065, w_005_066, w_005_067, w_005_068, w_005_069, w_005_070, w_005_071, w_005_072, w_005_073, w_005_074, w_005_075, w_005_076, w_005_077, w_005_078, w_005_080, w_005_081, w_005_082, w_005_083, w_005_084, w_005_085, w_005_086, w_005_087, w_005_088, w_005_089, w_005_090, w_005_091, w_005_092, w_005_093, w_005_094, w_005_095, w_005_096, w_005_097, w_005_098, w_005_099, w_005_100, w_005_101, w_005_103, w_005_104, w_005_105, w_005_106, w_005_107, w_005_108, w_005_109, w_005_110, w_005_111, w_005_112, w_005_113, w_005_114, w_005_115, w_005_117, w_005_118, w_005_119, w_005_120, w_005_121, w_005_122, w_005_123, w_005_124, w_005_125, w_005_126, w_005_127, w_005_130, w_005_132, w_005_133, w_005_134, w_005_135, w_005_136, w_005_137, w_005_138, w_005_139, w_005_141, w_005_142, w_005_143, w_005_144, w_005_145, w_005_146, w_005_147, w_005_148, w_005_149, w_005_150, w_005_151, w_005_152, w_005_153, w_005_154, w_005_155, w_005_156, w_005_157, w_005_158, w_005_159, w_005_160, w_005_161, w_005_162, w_005_163, w_005_164, w_005_165, w_005_166, w_005_167, w_005_168, w_005_169, w_005_170, w_005_171, w_005_172, w_005_173, w_005_175, w_005_176, w_005_177, w_005_178, w_005_179, w_005_180, w_005_181, w_005_182, w_005_184, w_005_185, w_005_186, w_005_187, w_005_188, w_005_189, w_005_190, w_005_191, w_005_192, w_005_193, w_005_194, w_005_195, w_005_196, w_005_197, w_005_198, w_005_199, w_005_200, w_005_201, w_005_203, w_005_206, w_005_207, w_005_208, w_005_210, w_005_211, w_005_212, w_005_213, w_005_214, w_005_215, w_005_216, w_005_217, w_005_218, w_005_219, w_005_220, w_005_221, w_005_222, w_005_223, w_005_224, w_005_225, w_005_226, w_005_227, w_005_228, w_005_229, w_005_230, w_005_231, w_005_232, w_005_233, w_005_235, w_005_236, w_005_237, w_005_238, w_005_239, w_005_241, w_005_242, w_005_243, w_005_244, w_005_245, w_005_246, w_005_250, w_005_251, w_005_252;
  wire w_006_000;
  wire w_007_001, w_007_002, w_007_003, w_007_004, w_007_005, w_007_006, w_007_007, w_007_008, w_007_009, w_007_013, w_007_014, w_007_015, w_007_016, w_007_017, w_007_018, w_007_019, w_007_020, w_007_021, w_007_022, w_007_023, w_007_025, w_007_026, w_007_027, w_007_029, w_007_030, w_007_031, w_007_032, w_007_033, w_007_035, w_007_038, w_007_039, w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045, w_007_046, w_007_047, w_007_048, w_007_049, w_007_050, w_007_051, w_007_052, w_007_053, w_007_055, w_007_056, w_007_057, w_007_058, w_007_059, w_007_060, w_007_061, w_007_062, w_007_063, w_007_064, w_007_065, w_007_066, w_007_068, w_007_069, w_007_070, w_007_071, w_007_072, w_007_073, w_007_074, w_007_075, w_007_076, w_007_077, w_007_078, w_007_080, w_007_081, w_007_082, w_007_083, w_007_084, w_007_085, w_007_086, w_007_087, w_007_088, w_007_089, w_007_090, w_007_091, w_007_092, w_007_094, w_007_095, w_007_097, w_007_098, w_007_099, w_007_100, w_007_101, w_007_104, w_007_105, w_007_106, w_007_107, w_007_108, w_007_109, w_007_113, w_007_115, w_007_116, w_007_117, w_007_118, w_007_119, w_007_120, w_007_121, w_007_122, w_007_123, w_007_124, w_007_125, w_007_126, w_007_128, w_007_129, w_007_131, w_007_134, w_007_135, w_007_136, w_007_137, w_007_138, w_007_141, w_007_142, w_007_143, w_007_144, w_007_146, w_007_147, w_007_148, w_007_154, w_007_156, w_007_159, w_007_160, w_007_163, w_007_164, w_007_165, w_007_166, w_007_167, w_007_168, w_007_170, w_007_171, w_007_172, w_007_173, w_007_174, w_007_175, w_007_176, w_007_177, w_007_178, w_007_180, w_007_181, w_007_182, w_007_183, w_007_184, w_007_186, w_007_187, w_007_188, w_007_189, w_007_190, w_007_192, w_007_193, w_007_194, w_007_195, w_007_196, w_007_197, w_007_199, w_007_200, w_007_203, w_007_204, w_007_206, w_007_208, w_007_209, w_007_210, w_007_211, w_007_213, w_007_214, w_007_215, w_007_216, w_007_219, w_007_221, w_007_222, w_007_224, w_007_225, w_007_226, w_007_227, w_007_228, w_007_229, w_007_230, w_007_231, w_007_233, w_007_234, w_007_238, w_007_239, w_007_240, w_007_241, w_007_242, w_007_243, w_007_244, w_007_245, w_007_246, w_007_247, w_007_248, w_007_249, w_007_250, w_007_251, w_007_252, w_007_253, w_007_254, w_007_255, w_007_258, w_007_259, w_007_260, w_007_261, w_007_262, w_007_263, w_007_264, w_007_265, w_007_266, w_007_267, w_007_268, w_007_269, w_007_270, w_007_271, w_007_272, w_007_273, w_007_275, w_007_276, w_007_278, w_007_281, w_007_283, w_007_284, w_007_285, w_007_286, w_007_288, w_007_290, w_007_292, w_007_293, w_007_296, w_007_297, w_007_298, w_007_299, w_007_300, w_007_302, w_007_303, w_007_305, w_007_306, w_007_307, w_007_308, w_007_309, w_007_314, w_007_315, w_007_316, w_007_317, w_007_319, w_007_320, w_007_321, w_007_322, w_007_324, w_007_325, w_007_328, w_007_329, w_007_333, w_007_337, w_007_340, w_007_341, w_007_342, w_007_343, w_007_344, w_007_345, w_007_347, w_007_348, w_007_349, w_007_350, w_007_352, w_007_354, w_007_355, w_007_356, w_007_357, w_007_359, w_007_360, w_007_361, w_007_362, w_007_363, w_007_364, w_007_366, w_007_367, w_007_368, w_007_370, w_007_371, w_007_372, w_007_373, w_007_374, w_007_376, w_007_377, w_007_378, w_007_379, w_007_380, w_007_381, w_007_382, w_007_383, w_007_385, w_007_386, w_007_388, w_007_389, w_007_390, w_007_391, w_007_394, w_007_396, w_007_398, w_007_400, w_007_403, w_007_404;
  wire w_008_000, w_008_001, w_008_003, w_008_004, w_008_005, w_008_008, w_008_010, w_008_011, w_008_012, w_008_013, w_008_014, w_008_015, w_008_016, w_008_017, w_008_018, w_008_020, w_008_022, w_008_023, w_008_024, w_008_025, w_008_026, w_008_027, w_008_028, w_008_029, w_008_030, w_008_031, w_008_032, w_008_033, w_008_034, w_008_035, w_008_037, w_008_038, w_008_039, w_008_040, w_008_041, w_008_043, w_008_045, w_008_046, w_008_047, w_008_048, w_008_050, w_008_051, w_008_052, w_008_053, w_008_054, w_008_056, w_008_057, w_008_058, w_008_059, w_008_060, w_008_061, w_008_062, w_008_063, w_008_064, w_008_065, w_008_066, w_008_067, w_008_068, w_008_070, w_008_072, w_008_073, w_008_074, w_008_075, w_008_076, w_008_077, w_008_078, w_008_079, w_008_080, w_008_081, w_008_082, w_008_083, w_008_084, w_008_085, w_008_086, w_008_087, w_008_088, w_008_089, w_008_090, w_008_091, w_008_092, w_008_093, w_008_095, w_008_096, w_008_098, w_008_099, w_008_100, w_008_102, w_008_103, w_008_104, w_008_105, w_008_106, w_008_107, w_008_109, w_008_110, w_008_111, w_008_112, w_008_113, w_008_114, w_008_115, w_008_116, w_008_117, w_008_118, w_008_119, w_008_120, w_008_121, w_008_123, w_008_124, w_008_125, w_008_126, w_008_127, w_008_128, w_008_130, w_008_131, w_008_132, w_008_133, w_008_134, w_008_135, w_008_137, w_008_138, w_008_139, w_008_140, w_008_142, w_008_143, w_008_145, w_008_146, w_008_148, w_008_149, w_008_150, w_008_152, w_008_153, w_008_154, w_008_156, w_008_157, w_008_161, w_008_162, w_008_165, w_008_166, w_008_168, w_008_169, w_008_173, w_008_175, w_008_176, w_008_177, w_008_179, w_008_180, w_008_183, w_008_184, w_008_185, w_008_186, w_008_187, w_008_190, w_008_191, w_008_193, w_008_195, w_008_196, w_008_198, w_008_199, w_008_200, w_008_201, w_008_202, w_008_203, w_008_205, w_008_206, w_008_207, w_008_208, w_008_209, w_008_210, w_008_212, w_008_215, w_008_216, w_008_218, w_008_219, w_008_223, w_008_225, w_008_226, w_008_228, w_008_230, w_008_231, w_008_233, w_008_234, w_008_236, w_008_237, w_008_238, w_008_239, w_008_240, w_008_241, w_008_242, w_008_243, w_008_244, w_008_245, w_008_246, w_008_250, w_008_251, w_008_252, w_008_253, w_008_254, w_008_255, w_008_256, w_008_258, w_008_260, w_008_261, w_008_263, w_008_264, w_008_268, w_008_269, w_008_270, w_008_271, w_008_273, w_008_274, w_008_275, w_008_276, w_008_277, w_008_280, w_008_282, w_008_283, w_008_287, w_008_288, w_008_290, w_008_291, w_008_292, w_008_294, w_008_296, w_008_297, w_008_299, w_008_300, w_008_302, w_008_304, w_008_307, w_008_309, w_008_310, w_008_311, w_008_312, w_008_315, w_008_317, w_008_318, w_008_320, w_008_321, w_008_324, w_008_325, w_008_327, w_008_329, w_008_331, w_008_333, w_008_337, w_008_342, w_008_343, w_008_345;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_004, w_009_005, w_009_006, w_009_007, w_009_008, w_009_009, w_009_010, w_009_011, w_009_012, w_009_013, w_009_014, w_009_015, w_009_016, w_009_017, w_009_018, w_009_019, w_009_020, w_009_021, w_009_022, w_009_024, w_009_025, w_009_026, w_009_027, w_009_028, w_009_029, w_009_030, w_009_031, w_009_032, w_009_033, w_009_034, w_009_035, w_009_036, w_009_037, w_009_038, w_009_040, w_009_041, w_009_042, w_009_043, w_009_044, w_009_045, w_009_046, w_009_047, w_009_048, w_009_049, w_009_050, w_009_051, w_009_052, w_009_054, w_009_056, w_009_058, w_009_059, w_009_061, w_009_062, w_009_063, w_009_064, w_009_065, w_009_067, w_009_072, w_009_073, w_009_074, w_009_075, w_009_076, w_009_077, w_009_078, w_009_079, w_009_080, w_009_081, w_009_083, w_009_084, w_009_086, w_009_088, w_009_089, w_009_090, w_009_091, w_009_092, w_009_093, w_009_094, w_009_096, w_009_098, w_009_099, w_009_101, w_009_103, w_009_104, w_009_105, w_009_106, w_009_107, w_009_108, w_009_109, w_009_111, w_009_112, w_009_113, w_009_115, w_009_116, w_009_117, w_009_118, w_009_120, w_009_121, w_009_122, w_009_123, w_009_124, w_009_125, w_009_126, w_009_127, w_009_128, w_009_129, w_009_130, w_009_131, w_009_132, w_009_133, w_009_134, w_009_135, w_009_136, w_009_137, w_009_139, w_009_140, w_009_142, w_009_143, w_009_144, w_009_145, w_009_146, w_009_147, w_009_148, w_009_149, w_009_151, w_009_152, w_009_153, w_009_154, w_009_155, w_009_156, w_009_157, w_009_158, w_009_159, w_009_160, w_009_161, w_009_162, w_009_163, w_009_164, w_009_165, w_009_167, w_009_168, w_009_169, w_009_170, w_009_171, w_009_172, w_009_173, w_009_174, w_009_175, w_009_176, w_009_177, w_009_178, w_009_179, w_009_181, w_009_183, w_009_185, w_009_186, w_009_187, w_009_189, w_009_190, w_009_191, w_009_192, w_009_193, w_009_194, w_009_196, w_009_197, w_009_198, w_009_199, w_009_200, w_009_202, w_009_203, w_009_204, w_009_206, w_009_208, w_009_209, w_009_211, w_009_212, w_009_213, w_009_216, w_009_217, w_009_218, w_009_220, w_009_221, w_009_222, w_009_223, w_009_224, w_009_225, w_009_226, w_009_227, w_009_228, w_009_229, w_009_231, w_009_232, w_009_233, w_009_234, w_009_235, w_009_236, w_009_237;
  wire w_010_002, w_010_004, w_010_005, w_010_007, w_010_008, w_010_009, w_010_012, w_010_013, w_010_014, w_010_015, w_010_016, w_010_018, w_010_020, w_010_021, w_010_023, w_010_024, w_010_025, w_010_026, w_010_027, w_010_028, w_010_029, w_010_030, w_010_033, w_010_034, w_010_035, w_010_036, w_010_037, w_010_038, w_010_040, w_010_041, w_010_042, w_010_044, w_010_045, w_010_046, w_010_047, w_010_048, w_010_049, w_010_051, w_010_052, w_010_053, w_010_054, w_010_055, w_010_059, w_010_062, w_010_063, w_010_064, w_010_065, w_010_067, w_010_069, w_010_071, w_010_072, w_010_073, w_010_075, w_010_076, w_010_077, w_010_078, w_010_079, w_010_083, w_010_087, w_010_089, w_010_094, w_010_096, w_010_097, w_010_098, w_010_100, w_010_101, w_010_103, w_010_104, w_010_107, w_010_108, w_010_112, w_010_115, w_010_116, w_010_119, w_010_120, w_010_121, w_010_123, w_010_127, w_010_128, w_010_131, w_010_132, w_010_134, w_010_135, w_010_136, w_010_137, w_010_142, w_010_144, w_010_145, w_010_146, w_010_150, w_010_151, w_010_152, w_010_153, w_010_158, w_010_159, w_010_162, w_010_163, w_010_170, w_010_172, w_010_174, w_010_175, w_010_176, w_010_178, w_010_179, w_010_180, w_010_181, w_010_185, w_010_187, w_010_188, w_010_189, w_010_190, w_010_191, w_010_192, w_010_193, w_010_196, w_010_197, w_010_198, w_010_201, w_010_204, w_010_207, w_010_208, w_010_211, w_010_213, w_010_214, w_010_216, w_010_217, w_010_218, w_010_219, w_010_220, w_010_223, w_010_224, w_010_225, w_010_226, w_010_234, w_010_235, w_010_236, w_010_240, w_010_241, w_010_244, w_010_246, w_010_247, w_010_251, w_010_253, w_010_254, w_010_255, w_010_256, w_010_258, w_010_260, w_010_261, w_010_262, w_010_263, w_010_264, w_010_265, w_010_266, w_010_267, w_010_268, w_010_270, w_010_273, w_010_276, w_010_278, w_010_281, w_010_282, w_010_283, w_010_284, w_010_286, w_010_287, w_010_288, w_010_289, w_010_290, w_010_291, w_010_292, w_010_294, w_010_298, w_010_303, w_010_304, w_010_306, w_010_307, w_010_309, w_010_311, w_010_315, w_010_316, w_010_317, w_010_318, w_010_321, w_010_322, w_010_323, w_010_325, w_010_326, w_010_327, w_010_328, w_010_332, w_010_333, w_010_334, w_010_336, w_010_337, w_010_338, w_010_342, w_010_343, w_010_344, w_010_345, w_010_346, w_010_347, w_010_348, w_010_349, w_010_351, w_010_353, w_010_354, w_010_357, w_010_359, w_010_361, w_010_362, w_010_364, w_010_368, w_010_372, w_010_377, w_010_379, w_010_380, w_010_381, w_010_382, w_010_384, w_010_385, w_010_389, w_010_391, w_010_392, w_010_398, w_010_400, w_010_402, w_010_404, w_010_406, w_010_408, w_010_410, w_010_412, w_010_413, w_010_416, w_010_417, w_010_418, w_010_422, w_010_423, w_010_425, w_010_427, w_010_429, w_010_431, w_010_433, w_010_435, w_010_436, w_010_438, w_010_441, w_010_443, w_010_445, w_010_446, w_010_448, w_010_449, w_010_450, w_010_451;
  wire w_011_000, w_011_001, w_011_004, w_011_009, w_011_011, w_011_012, w_011_014, w_011_015, w_011_016, w_011_017, w_011_018, w_011_019, w_011_020, w_011_021, w_011_022, w_011_023, w_011_025, w_011_026, w_011_027, w_011_028, w_011_030, w_011_031, w_011_033, w_011_034, w_011_035, w_011_036, w_011_037, w_011_038, w_011_039, w_011_041, w_011_042, w_011_043, w_011_045, w_011_047, w_011_051, w_011_052, w_011_053, w_011_054, w_011_055, w_011_056, w_011_057, w_011_058, w_011_059, w_011_060, w_011_061, w_011_063, w_011_064, w_011_066, w_011_067, w_011_068, w_011_069, w_011_071, w_011_072, w_011_073, w_011_076, w_011_077, w_011_078, w_011_079, w_011_080, w_011_081, w_011_082, w_011_083, w_011_084, w_011_085, w_011_086, w_011_087, w_011_088, w_011_089, w_011_090, w_011_091, w_011_092, w_011_093, w_011_095, w_011_096, w_011_097, w_011_098, w_011_099, w_011_100, w_011_101, w_011_102, w_011_104, w_011_106, w_011_108, w_011_110, w_011_111, w_011_112, w_011_113, w_011_114, w_011_115, w_011_116, w_011_117, w_011_120, w_011_121, w_011_123, w_011_124, w_011_125, w_011_126, w_011_127, w_011_128, w_011_130, w_011_131, w_011_132, w_011_133, w_011_134, w_011_135, w_011_136, w_011_137, w_011_140, w_011_141, w_011_142, w_011_143, w_011_144, w_011_146, w_011_150, w_011_151, w_011_152, w_011_153, w_011_155, w_011_156, w_011_159, w_011_160, w_011_161, w_011_163, w_011_164, w_011_166, w_011_169, w_011_177, w_011_178, w_011_179, w_011_181, w_011_182, w_011_183, w_011_186, w_011_187, w_011_188, w_011_189, w_011_192, w_011_194, w_011_196, w_011_197, w_011_200, w_011_201, w_011_204, w_011_205, w_011_206, w_011_207, w_011_211, w_011_213, w_011_214, w_011_215, w_011_218, w_011_219, w_011_220, w_011_221, w_011_222, w_011_224, w_011_226, w_011_228, w_011_230, w_011_231, w_011_232, w_011_233, w_011_234, w_011_238, w_011_242, w_011_246, w_011_249, w_011_251, w_011_253, w_011_254, w_011_257, w_011_268, w_011_269, w_011_272, w_011_273, w_011_276, w_011_278, w_011_279, w_011_280, w_011_282, w_011_284, w_011_285, w_011_286, w_011_287, w_011_289, w_011_291, w_011_292, w_011_294, w_011_295, w_011_296, w_011_297, w_011_300, w_011_301, w_011_303, w_011_304, w_011_308, w_011_309, w_011_312, w_011_315, w_011_317, w_011_318, w_011_319, w_011_320, w_011_321, w_011_323, w_011_327, w_011_329, w_011_331, w_011_332, w_011_333, w_011_334, w_011_335, w_011_336, w_011_337, w_011_339, w_011_340, w_011_342;
  wire w_012_000, w_012_001, w_012_002, w_012_003, w_012_004, w_012_005, w_012_006, w_012_007, w_012_010, w_012_012, w_012_013, w_012_014, w_012_015, w_012_016, w_012_017, w_012_018, w_012_019, w_012_020, w_012_021, w_012_023, w_012_024, w_012_025, w_012_026, w_012_027, w_012_028, w_012_029, w_012_030, w_012_031, w_012_032, w_012_034, w_012_035, w_012_036, w_012_038, w_012_039, w_012_040, w_012_041, w_012_042, w_012_043, w_012_045, w_012_046, w_012_048, w_012_049, w_012_050, w_012_052, w_012_053, w_012_054, w_012_055, w_012_056, w_012_057, w_012_060, w_012_061, w_012_063, w_012_065, w_012_067, w_012_068, w_012_070, w_012_071, w_012_073, w_012_074, w_012_077, w_012_080, w_012_081, w_012_083, w_012_084, w_012_086, w_012_088, w_012_089, w_012_090, w_012_091, w_012_092, w_012_094, w_012_096, w_012_097, w_012_098, w_012_099, w_012_101, w_012_103, w_012_108, w_012_109, w_012_110, w_012_113, w_012_114, w_012_116, w_012_119, w_012_122, w_012_125, w_012_126, w_012_127, w_012_131, w_012_132, w_012_133, w_012_135, w_012_138, w_012_143, w_012_144, w_012_146, w_012_147, w_012_149, w_012_151, w_012_158, w_012_159, w_012_160, w_012_161, w_012_165, w_012_166, w_012_169, w_012_170, w_012_171, w_012_174, w_012_175, w_012_176, w_012_177, w_012_178, w_012_180, w_012_181, w_012_182, w_012_184, w_012_186, w_012_187, w_012_189, w_012_191, w_012_195, w_012_197, w_012_200, w_012_201, w_012_205, w_012_211, w_012_212, w_012_214, w_012_215, w_012_217, w_012_218, w_012_219, w_012_220, w_012_221, w_012_222, w_012_223, w_012_225, w_012_226, w_012_227, w_012_230, w_012_234, w_012_236, w_012_238, w_012_239, w_012_241, w_012_245, w_012_248, w_012_249, w_012_250, w_012_253, w_012_255, w_012_256, w_012_258, w_012_260, w_012_261, w_012_262, w_012_263, w_012_265, w_012_266, w_012_270, w_012_272, w_012_275, w_012_277, w_012_278, w_012_279, w_012_280, w_012_282, w_012_283, w_012_284, w_012_285, w_012_286, w_012_290, w_012_291, w_012_293, w_012_294, w_012_295, w_012_296, w_012_298, w_012_300, w_012_303, w_012_309, w_012_310, w_012_312, w_012_313, w_012_314, w_012_315, w_012_318, w_012_320, w_012_321, w_012_322, w_012_324, w_012_325, w_012_326, w_012_328, w_012_330, w_012_333, w_012_336, w_012_337, w_012_339, w_012_340, w_012_341, w_012_344, w_012_345, w_012_347, w_012_348, w_012_349, w_012_350, w_012_353, w_012_356, w_012_357, w_012_358, w_012_359, w_012_362, w_012_363, w_012_364, w_012_365, w_012_366, w_012_367, w_012_368, w_012_369, w_012_373, w_012_374, w_012_379, w_012_380, w_012_382;
  wire w_013_000, w_013_001, w_013_005, w_013_006, w_013_007, w_013_008, w_013_009, w_013_010, w_013_011, w_013_012, w_013_013, w_013_014, w_013_017, w_013_018, w_013_019, w_013_020, w_013_022, w_013_023, w_013_024, w_013_025, w_013_027, w_013_028, w_013_030, w_013_032, w_013_033, w_013_034, w_013_035, w_013_036, w_013_037, w_013_038, w_013_039, w_013_040, w_013_041, w_013_043, w_013_044, w_013_046, w_013_047, w_013_049, w_013_050, w_013_051, w_013_052, w_013_053, w_013_054, w_013_055, w_013_057, w_013_059, w_013_060, w_013_061, w_013_062, w_013_063, w_013_065, w_013_066, w_013_068, w_013_071, w_013_073, w_013_075, w_013_080, w_013_081, w_013_082, w_013_083, w_013_084, w_013_087, w_013_088, w_013_089, w_013_090, w_013_091, w_013_093, w_013_094, w_013_095, w_013_096, w_013_097, w_013_099, w_013_100, w_013_101, w_013_102, w_013_103, w_013_104, w_013_105, w_013_106, w_013_108, w_013_109, w_013_110, w_013_112, w_013_113, w_013_116, w_013_117, w_013_118, w_013_119, w_013_120, w_013_122, w_013_123, w_013_124, w_013_126, w_013_127, w_013_129, w_013_132, w_013_133, w_013_134, w_013_135, w_013_140, w_013_141, w_013_142, w_013_144, w_013_145, w_013_146, w_013_147, w_013_148, w_013_149, w_013_150, w_013_151, w_013_152, w_013_153, w_013_154, w_013_155, w_013_158, w_013_159, w_013_160, w_013_161, w_013_162, w_013_163, w_013_164, w_013_165, w_013_166, w_013_167, w_013_168, w_013_169, w_013_171, w_013_172, w_013_173, w_013_174, w_013_175, w_013_176, w_013_177, w_013_180, w_013_181, w_013_182, w_013_183, w_013_184, w_013_185, w_013_186, w_013_187, w_013_188, w_013_189, w_013_190, w_013_191, w_013_192, w_013_193, w_013_194, w_013_195, w_013_196, w_013_197, w_013_199, w_013_200, w_013_201, w_013_204, w_013_205, w_013_207, w_013_208, w_013_210, w_013_211, w_013_213, w_013_214, w_013_215, w_013_217, w_013_218, w_013_220, w_013_221, w_013_222, w_013_223, w_013_224, w_013_225, w_013_226, w_013_227, w_013_228, w_013_229, w_013_231, w_013_232, w_013_235, w_013_239, w_013_243, w_013_245, w_013_246, w_013_248, w_013_250, w_013_253, w_013_255, w_013_261, w_013_264, w_013_265, w_013_266, w_013_267, w_013_268;
  wire w_014_001, w_014_002, w_014_005, w_014_006, w_014_007, w_014_008, w_014_009, w_014_010, w_014_011, w_014_013, w_014_014, w_014_016, w_014_017, w_014_018, w_014_020, w_014_022, w_014_023, w_014_024, w_014_025, w_014_027, w_014_028, w_014_033, w_014_034, w_014_035, w_014_037, w_014_038, w_014_039, w_014_040, w_014_043, w_014_044, w_014_045, w_014_046, w_014_047, w_014_048, w_014_049, w_014_052, w_014_053, w_014_054, w_014_056, w_014_057, w_014_058, w_014_059, w_014_060, w_014_063, w_014_065, w_014_066, w_014_067, w_014_068, w_014_069, w_014_070, w_014_071, w_014_072, w_014_073, w_014_074, w_014_076, w_014_079, w_014_080, w_014_081, w_014_082, w_014_083, w_014_084, w_014_085, w_014_086, w_014_087, w_014_088, w_014_091, w_014_092, w_014_093, w_014_094, w_014_095, w_014_096, w_014_099, w_014_101, w_014_102, w_014_103, w_014_104, w_014_105, w_014_106, w_014_108, w_014_109, w_014_110, w_014_113, w_014_114, w_014_115, w_014_116, w_014_118, w_014_119, w_014_121, w_014_122, w_014_123, w_014_125, w_014_128, w_014_129, w_014_131, w_014_132, w_014_133, w_014_134, w_014_135, w_014_136, w_014_137, w_014_138, w_014_140, w_014_141, w_014_144, w_014_145, w_014_146, w_014_148, w_014_150, w_014_151, w_014_152, w_014_153, w_014_154, w_014_155, w_014_156, w_014_157, w_014_159, w_014_161, w_014_163, w_014_164, w_014_165, w_014_166, w_014_167, w_014_169, w_014_170, w_014_173, w_014_174, w_014_178, w_014_181, w_014_182, w_014_183, w_014_184, w_014_185, w_014_186, w_014_188, w_014_191, w_014_193, w_014_195, w_014_196, w_014_197, w_014_198, w_014_202, w_014_203, w_014_204, w_014_205, w_014_206, w_014_207, w_014_208, w_014_209, w_014_210, w_014_211, w_014_212, w_014_213, w_014_215, w_014_216, w_014_217, w_014_218, w_014_219, w_014_220, w_014_221, w_014_222, w_014_225, w_014_226, w_014_227, w_014_228, w_014_229, w_014_231, w_014_233, w_014_234, w_014_235, w_014_236, w_014_237, w_014_240, w_014_241, w_014_243, w_014_245, w_014_247, w_014_248, w_014_249, w_014_252, w_014_254, w_014_256, w_014_259, w_014_260, w_014_262, w_014_264, w_014_265;
  wire w_015_000, w_015_001, w_015_002, w_015_004, w_015_005, w_015_006, w_015_007, w_015_009, w_015_010, w_015_011, w_015_012, w_015_013, w_015_014, w_015_015, w_015_017, w_015_018, w_015_020, w_015_021, w_015_022, w_015_023, w_015_024, w_015_025, w_015_026, w_015_027, w_015_028, w_015_029, w_015_031, w_015_033, w_015_034, w_015_036, w_015_037, w_015_038, w_015_039, w_015_040, w_015_041, w_015_042, w_015_043, w_015_044, w_015_045, w_015_046, w_015_047, w_015_048, w_015_049, w_015_050, w_015_051, w_015_052, w_015_053, w_015_054, w_015_055, w_015_058, w_015_059, w_015_060, w_015_061, w_015_062, w_015_063, w_015_064, w_015_065, w_015_066, w_015_067, w_015_068, w_015_069, w_015_070, w_015_071, w_015_072, w_015_073, w_015_074, w_015_075, w_015_077, w_015_078, w_015_080, w_015_081, w_015_082, w_015_083, w_015_085, w_015_086, w_015_088, w_015_089, w_015_090, w_015_091, w_015_092, w_015_093, w_015_095, w_015_096, w_015_097, w_015_098, w_015_100, w_015_102, w_015_105, w_015_106, w_015_108, w_015_111, w_015_112, w_015_113, w_015_114, w_015_115, w_015_116, w_015_117, w_015_120, w_015_121, w_015_122, w_015_124, w_015_125, w_015_126, w_015_127, w_015_128, w_015_129, w_015_131, w_015_132, w_015_134;
  wire w_016_001, w_016_002, w_016_003, w_016_005, w_016_007, w_016_008, w_016_009, w_016_011, w_016_012, w_016_014, w_016_015, w_016_016, w_016_017, w_016_018, w_016_019, w_016_020, w_016_021, w_016_022, w_016_023, w_016_024, w_016_026, w_016_027, w_016_028, w_016_029, w_016_030, w_016_031, w_016_032, w_016_033, w_016_034, w_016_035, w_016_037, w_016_038, w_016_044, w_016_045, w_016_046, w_016_048, w_016_049, w_016_051, w_016_052, w_016_053, w_016_056, w_016_058, w_016_059, w_016_061, w_016_062, w_016_065, w_016_067, w_016_068, w_016_070, w_016_071, w_016_073, w_016_074, w_016_076, w_016_077, w_016_078, w_016_079, w_016_080, w_016_082, w_016_084, w_016_085, w_016_086, w_016_087, w_016_091, w_016_093, w_016_094, w_016_095, w_016_097, w_016_099, w_016_101, w_016_106, w_016_107, w_016_110, w_016_111, w_016_113, w_016_117, w_016_118, w_016_119, w_016_122, w_016_124, w_016_125, w_016_130, w_016_133, w_016_136, w_016_139, w_016_140, w_016_141, w_016_144, w_016_145, w_016_147, w_016_149, w_016_151, w_016_152, w_016_153, w_016_157, w_016_164, w_016_165, w_016_169, w_016_173, w_016_175, w_016_176, w_016_177, w_016_178, w_016_182, w_016_183, w_016_185, w_016_187, w_016_189, w_016_191, w_016_192, w_016_194, w_016_197, w_016_200, w_016_209, w_016_210, w_016_212, w_016_213, w_016_214, w_016_216, w_016_222, w_016_223, w_016_225, w_016_228, w_016_230, w_016_232, w_016_233, w_016_234, w_016_239, w_016_241, w_016_244, w_016_245, w_016_247, w_016_248, w_016_249, w_016_250, w_016_253, w_016_254, w_016_255, w_016_256, w_016_257, w_016_258, w_016_260, w_016_262, w_016_263, w_016_264, w_016_265, w_016_268, w_016_274, w_016_278, w_016_279, w_016_280, w_016_281, w_016_285, w_016_286, w_016_287, w_016_291, w_016_292, w_016_294, w_016_295, w_016_297, w_016_300, w_016_301, w_016_303, w_016_304, w_016_310, w_016_311, w_016_315, w_016_316, w_016_319, w_016_322, w_016_324, w_016_328, w_016_330, w_016_335, w_016_336, w_016_337, w_016_339, w_016_345, w_016_347, w_016_349, w_016_350, w_016_354, w_016_355, w_016_356, w_016_357, w_016_362, w_016_364, w_016_367, w_016_369, w_016_371, w_016_372, w_016_374, w_016_375, w_016_378, w_016_380, w_016_381, w_016_382, w_016_384, w_016_385, w_016_391, w_016_394, w_016_395, w_016_398, w_016_399;
  wire w_017_000, w_017_001, w_017_003, w_017_004, w_017_005, w_017_006, w_017_007, w_017_008, w_017_009, w_017_010, w_017_011, w_017_012, w_017_014, w_017_015, w_017_016, w_017_017, w_017_018, w_017_019, w_017_020, w_017_021, w_017_022, w_017_023, w_017_024, w_017_025, w_017_026, w_017_027, w_017_028, w_017_029, w_017_030, w_017_033, w_017_034, w_017_035, w_017_036, w_017_037, w_017_038, w_017_039, w_017_040, w_017_041, w_017_042, w_017_043, w_017_044, w_017_045, w_017_046, w_017_047, w_017_048, w_017_049, w_017_050, w_017_051, w_017_052, w_017_053, w_017_054, w_017_055, w_017_056, w_017_058, w_017_059, w_017_060, w_017_061, w_017_063, w_017_064, w_017_065, w_017_066, w_017_067, w_017_070, w_017_071, w_017_072, w_017_073, w_017_074, w_017_075, w_017_076, w_017_077, w_017_078, w_017_080, w_017_081, w_017_083, w_017_084, w_017_085, w_017_086, w_017_087, w_017_088, w_017_091, w_017_092, w_017_093, w_017_094, w_017_098, w_017_099, w_017_100, w_017_101, w_017_103, w_017_104, w_017_108, w_017_109, w_017_111, w_017_113, w_017_114, w_017_115, w_017_116, w_017_117, w_017_118, w_017_122, w_017_123, w_017_124, w_017_126, w_017_128, w_017_130, w_017_133, w_017_135, w_017_136, w_017_138, w_017_139, w_017_141, w_017_143, w_017_144, w_017_146, w_017_148, w_017_150, w_017_154, w_017_155, w_017_156, w_017_157, w_017_159, w_017_162, w_017_163, w_017_166, w_017_167, w_017_168, w_017_171, w_017_172, w_017_173, w_017_176, w_017_177, w_017_178, w_017_179, w_017_180, w_017_181, w_017_182, w_017_184, w_017_185, w_017_186, w_017_187, w_017_188, w_017_190, w_017_191;
  wire w_018_000, w_018_001, w_018_002, w_018_003, w_018_005, w_018_006, w_018_008, w_018_010, w_018_012, w_018_014, w_018_015, w_018_016, w_018_017, w_018_018, w_018_019, w_018_020, w_018_022, w_018_023, w_018_026, w_018_027, w_018_030, w_018_031, w_018_032, w_018_034, w_018_035, w_018_037, w_018_039, w_018_040, w_018_045, w_018_047, w_018_048, w_018_050, w_018_051, w_018_053, w_018_054, w_018_057, w_018_059, w_018_060, w_018_061, w_018_063, w_018_064, w_018_067, w_018_068, w_018_070, w_018_071, w_018_072, w_018_074, w_018_075, w_018_076, w_018_078, w_018_080, w_018_081, w_018_083, w_018_084, w_018_086, w_018_089, w_018_091, w_018_094, w_018_095, w_018_096, w_018_097, w_018_098, w_018_100, w_018_102, w_018_103, w_018_104, w_018_105, w_018_106, w_018_107, w_018_108, w_018_110, w_018_111, w_018_112, w_018_114, w_018_118, w_018_119, w_018_123, w_018_124, w_018_125, w_018_126, w_018_127, w_018_130, w_018_131, w_018_132, w_018_133, w_018_134, w_018_135, w_018_136, w_018_137, w_018_139, w_018_141, w_018_142, w_018_143, w_018_144, w_018_145, w_018_146, w_018_150, w_018_151, w_018_153, w_018_155, w_018_156, w_018_157, w_018_158, w_018_160, w_018_161, w_018_162, w_018_163, w_018_164, w_018_165, w_018_167, w_018_168, w_018_169, w_018_171, w_018_173, w_018_175, w_018_181, w_018_182, w_018_183, w_018_186, w_018_187, w_018_196, w_018_197, w_018_199, w_018_200, w_018_203, w_018_206, w_018_211, w_018_212, w_018_213, w_018_215, w_018_218, w_018_229, w_018_234, w_018_235, w_018_236, w_018_237, w_018_239, w_018_243, w_018_246, w_018_248, w_018_249, w_018_250, w_018_256, w_018_257, w_018_259, w_018_263, w_018_270, w_018_278, w_018_279, w_018_282, w_018_283, w_018_285, w_018_287, w_018_288, w_018_291, w_018_292, w_018_293, w_018_295, w_018_297, w_018_300, w_018_301, w_018_302, w_018_306, w_018_311, w_018_312, w_018_313, w_018_314, w_018_320, w_018_321, w_018_322;
  wire w_019_000, w_019_001, w_019_002, w_019_003, w_019_004, w_019_005, w_019_006, w_019_007, w_019_008, w_019_009, w_019_010, w_019_011, w_019_012, w_019_013, w_019_014, w_019_015, w_019_016, w_019_017, w_019_018, w_019_019, w_019_020, w_019_021, w_019_022, w_019_023, w_019_024, w_019_025, w_019_026, w_019_027, w_019_028, w_019_029, w_019_030, w_019_031, w_019_032, w_019_033, w_019_034, w_019_035, w_019_036, w_019_037, w_019_038, w_019_039, w_019_040, w_019_041, w_019_042, w_019_043, w_019_044, w_019_045, w_019_046, w_019_047, w_019_048, w_019_049, w_019_050, w_019_051, w_019_052, w_019_053;
  wire w_020_000, w_020_001, w_020_003, w_020_005, w_020_007, w_020_009, w_020_011, w_020_012, w_020_013, w_020_014, w_020_015, w_020_016, w_020_019, w_020_020, w_020_022, w_020_023, w_020_024, w_020_025, w_020_026, w_020_028, w_020_030, w_020_031, w_020_032, w_020_033, w_020_034, w_020_035, w_020_037, w_020_038, w_020_039, w_020_040, w_020_042, w_020_043, w_020_044, w_020_045, w_020_046, w_020_048, w_020_049, w_020_050, w_020_051, w_020_052, w_020_053, w_020_054, w_020_055, w_020_056, w_020_059, w_020_060, w_020_062, w_020_063, w_020_065, w_020_066, w_020_068, w_020_069, w_020_071, w_020_072, w_020_073, w_020_074, w_020_075, w_020_078, w_020_079, w_020_080, w_020_083, w_020_084, w_020_085, w_020_086, w_020_088, w_020_089, w_020_091, w_020_094, w_020_095, w_020_096, w_020_097, w_020_098, w_020_099, w_020_100, w_020_101, w_020_103, w_020_104, w_020_105, w_020_106, w_020_107, w_020_108, w_020_112, w_020_113, w_020_114, w_020_115, w_020_117, w_020_119, w_020_120, w_020_123, w_020_124, w_020_125, w_020_126, w_020_127, w_020_128, w_020_131, w_020_135, w_020_136, w_020_137, w_020_138, w_020_139, w_020_140, w_020_145, w_020_146, w_020_150, w_020_151, w_020_152, w_020_153, w_020_154, w_020_155, w_020_156, w_020_157, w_020_158, w_020_159, w_020_161, w_020_162, w_020_163, w_020_164, w_020_165, w_020_167, w_020_170, w_020_171, w_020_172, w_020_173, w_020_175, w_020_176, w_020_180, w_020_182, w_020_183, w_020_184, w_020_186;
  wire w_021_000, w_021_001, w_021_002, w_021_003, w_021_005, w_021_007, w_021_008, w_021_009, w_021_010, w_021_011, w_021_012, w_021_014, w_021_015, w_021_016, w_021_017, w_021_018, w_021_020, w_021_021, w_021_022, w_021_023, w_021_024, w_021_025, w_021_026, w_021_027, w_021_028, w_021_029, w_021_030, w_021_031, w_021_032, w_021_033, w_021_034, w_021_035, w_021_036, w_021_037, w_021_038, w_021_039, w_021_040, w_021_041, w_021_042, w_021_043, w_021_044, w_021_045, w_021_047, w_021_048, w_021_049, w_021_050, w_021_051, w_021_052, w_021_053, w_021_056, w_021_057, w_021_058, w_021_059, w_021_060, w_021_061, w_021_063, w_021_064, w_021_066, w_021_067, w_021_069, w_021_070, w_021_071, w_021_072, w_021_073, w_021_075, w_021_076, w_021_077, w_021_078, w_021_079, w_021_081, w_021_082, w_021_083, w_021_084, w_021_085, w_021_086, w_021_088, w_021_089, w_021_090, w_021_091, w_021_092, w_021_093, w_021_094, w_021_096, w_021_097, w_021_098, w_021_099, w_021_100, w_021_101, w_021_102, w_021_103, w_021_104, w_021_105, w_021_106, w_021_107, w_021_108, w_021_109;
  wire w_022_000, w_022_002, w_022_003, w_022_004, w_022_005, w_022_006, w_022_007, w_022_009, w_022_010, w_022_011, w_022_012, w_022_013, w_022_014, w_022_016, w_022_018, w_022_020, w_022_021, w_022_023, w_022_024, w_022_025, w_022_027, w_022_028, w_022_032, w_022_033, w_022_034, w_022_035, w_022_036, w_022_037, w_022_038, w_022_040, w_022_041, w_022_042, w_022_043, w_022_044, w_022_046, w_022_049, w_022_050, w_022_051, w_022_052, w_022_053, w_022_055, w_022_056, w_022_057, w_022_058, w_022_059, w_022_062, w_022_064, w_022_065, w_022_067, w_022_069, w_022_070, w_022_071, w_022_072, w_022_074, w_022_075, w_022_076, w_022_078, w_022_079, w_022_081, w_022_082, w_022_083, w_022_084, w_022_085, w_022_088, w_022_090, w_022_091, w_022_092, w_022_093, w_022_095, w_022_096, w_022_098, w_022_099, w_022_101, w_022_102, w_022_103, w_022_105, w_022_106, w_022_107, w_022_109, w_022_110, w_022_112, w_022_113, w_022_114, w_022_115, w_022_116, w_022_117, w_022_118, w_022_120, w_022_121, w_022_122, w_022_123, w_022_124, w_022_126, w_022_127, w_022_131, w_022_132, w_022_133, w_022_134, w_022_137, w_022_138, w_022_139, w_022_140, w_022_141, w_022_142, w_022_143, w_022_144, w_022_145, w_022_146, w_022_147, w_022_148, w_022_149, w_022_152, w_022_154, w_022_156, w_022_157, w_022_158, w_022_159, w_022_160, w_022_161, w_022_162, w_022_164, w_022_165, w_022_166, w_022_167, w_022_168, w_022_169, w_022_170, w_022_171, w_022_172, w_022_173;
  wire w_023_000, w_023_002, w_023_006, w_023_009, w_023_010, w_023_013, w_023_014, w_023_016, w_023_018, w_023_020, w_023_024, w_023_028, w_023_030, w_023_031, w_023_034, w_023_038, w_023_039, w_023_041, w_023_042, w_023_043, w_023_046, w_023_047, w_023_049, w_023_050, w_023_051, w_023_052, w_023_053, w_023_058, w_023_059, w_023_061, w_023_063, w_023_064, w_023_067, w_023_068, w_023_071, w_023_072, w_023_074, w_023_075, w_023_081, w_023_082, w_023_083, w_023_100, w_023_104, w_023_110, w_023_120, w_023_121, w_023_122, w_023_126, w_023_137, w_023_138, w_023_140, w_023_144, w_023_145, w_023_150, w_023_156, w_023_159, w_023_161, w_023_163, w_023_165, w_023_172, w_023_176, w_023_177, w_023_179, w_023_180, w_023_182, w_023_183, w_023_185, w_023_189, w_023_190, w_023_191, w_023_192, w_023_196, w_023_197, w_023_201, w_023_209, w_023_210, w_023_215, w_023_218, w_023_220, w_023_228, w_023_231, w_023_232, w_023_233, w_023_235, w_023_238, w_023_239, w_023_244, w_023_251, w_023_256, w_023_259, w_023_264, w_023_267, w_023_269, w_023_270, w_023_271, w_023_272, w_023_275, w_023_277, w_023_284, w_023_285, w_023_290, w_023_295, w_023_301, w_023_306, w_023_307, w_023_309, w_023_311, w_023_312, w_023_314, w_023_318, w_023_319, w_023_323, w_023_324, w_023_325, w_023_327, w_023_330, w_023_334, w_023_335, w_023_340, w_023_348, w_023_350, w_023_351, w_023_353, w_023_354, w_023_359, w_023_367, w_023_369, w_023_373, w_023_374, w_023_376, w_023_379, w_023_386, w_023_388, w_023_393, w_023_395, w_023_400, w_023_401, w_023_402, w_023_404, w_023_413;
  wire w_024_000, w_024_002, w_024_003, w_024_004, w_024_007, w_024_008, w_024_009, w_024_016, w_024_018, w_024_019, w_024_021, w_024_023, w_024_025, w_024_027, w_024_031, w_024_032, w_024_033, w_024_036, w_024_037, w_024_040, w_024_042, w_024_044, w_024_045, w_024_046, w_024_048, w_024_049, w_024_051, w_024_052, w_024_053, w_024_054, w_024_055, w_024_057, w_024_058, w_024_059, w_024_060, w_024_061, w_024_064, w_024_065, w_024_066, w_024_067, w_024_068, w_024_069, w_024_070, w_024_071, w_024_072, w_024_073, w_024_074, w_024_075, w_024_076, w_024_078, w_024_081, w_024_084, w_024_085, w_024_086, w_024_087, w_024_088, w_024_089, w_024_090, w_024_093, w_024_096, w_024_100, w_024_103, w_024_105, w_024_106, w_024_109, w_024_110, w_024_111, w_024_112, w_024_114, w_024_115, w_024_116, w_024_117, w_024_121, w_024_122, w_024_123, w_024_124, w_024_127, w_024_128, w_024_130, w_024_131, w_024_132, w_024_133, w_024_135, w_024_136, w_024_139, w_024_140, w_024_143, w_024_144, w_024_148, w_024_150, w_024_151, w_024_152, w_024_153, w_024_163, w_024_164, w_024_165, w_024_166, w_024_169, w_024_170, w_024_173, w_024_174, w_024_176, w_024_177, w_024_178, w_024_179, w_024_180, w_024_181, w_024_182, w_024_183, w_024_185, w_024_186, w_024_187, w_024_188, w_024_189, w_024_190, w_024_191, w_024_194, w_024_196, w_024_197, w_024_205, w_024_206, w_024_209, w_024_210, w_024_211, w_024_214, w_024_216, w_024_217, w_024_222, w_024_226, w_024_228, w_024_229, w_024_230, w_024_235, w_024_239, w_024_240, w_024_241, w_024_244, w_024_245, w_024_249, w_024_250, w_024_251, w_024_258, w_024_259, w_024_261, w_024_266, w_024_270, w_024_275, w_024_276, w_024_277, w_024_280, w_024_284, w_024_285, w_024_287, w_024_294, w_024_295, w_024_296, w_024_297;
  wire w_025_007, w_025_009, w_025_010, w_025_012, w_025_013, w_025_014, w_025_015, w_025_016, w_025_017, w_025_019, w_025_020, w_025_023, w_025_026, w_025_029, w_025_030, w_025_045, w_025_056, w_025_060, w_025_063, w_025_066, w_025_069, w_025_070, w_025_071, w_025_073, w_025_074, w_025_079, w_025_082, w_025_085, w_025_089, w_025_091, w_025_092, w_025_093, w_025_094, w_025_095, w_025_097, w_025_101, w_025_104, w_025_105, w_025_106, w_025_113, w_025_115, w_025_127, w_025_130, w_025_137, w_025_143, w_025_146, w_025_149, w_025_150, w_025_155, w_025_156, w_025_159, w_025_160, w_025_165, w_025_172, w_025_174, w_025_180, w_025_190, w_025_194, w_025_195, w_025_197, w_025_200, w_025_212, w_025_214, w_025_220, w_025_226, w_025_233, w_025_234, w_025_237, w_025_240, w_025_244, w_025_245, w_025_248, w_025_249, w_025_258, w_025_260, w_025_261, w_025_262, w_025_264, w_025_265, w_025_275, w_025_276, w_025_277, w_025_279, w_025_282, w_025_285, w_025_287, w_025_288, w_025_293, w_025_295, w_025_297, w_025_311, w_025_315, w_025_318, w_025_320, w_025_321, w_025_322, w_025_325, w_025_326, w_025_331, w_025_333, w_025_336, w_025_340, w_025_349, w_025_350, w_025_354, w_025_359, w_025_362, w_025_373, w_025_375, w_025_376, w_025_380, w_025_385, w_025_388, w_025_391, w_025_394, w_025_396, w_025_402, w_025_404, w_025_413, w_025_416, w_025_420, w_025_422, w_025_423, w_025_424, w_025_428, w_025_429, w_025_431, w_025_445, w_025_446, w_025_450, w_025_456, w_025_459, w_025_463, w_025_466, w_025_470, w_025_471, w_025_472, w_025_476, w_025_477;
  wire w_026_002, w_026_003, w_026_004, w_026_007, w_026_011, w_026_012, w_026_013, w_026_014, w_026_017, w_026_018, w_026_020, w_026_021, w_026_022, w_026_025, w_026_033, w_026_034, w_026_035, w_026_036, w_026_038, w_026_039, w_026_042, w_026_048, w_026_049, w_026_050, w_026_056, w_026_058, w_026_060, w_026_066, w_026_068, w_026_070, w_026_072, w_026_073, w_026_082, w_026_084, w_026_087, w_026_088, w_026_091, w_026_098, w_026_099, w_026_102, w_026_103, w_026_104, w_026_105, w_026_113, w_026_114, w_026_118, w_026_125, w_026_127, w_026_128, w_026_131, w_026_133, w_026_137, w_026_142, w_026_145, w_026_148, w_026_150, w_026_151, w_026_162, w_026_173, w_026_175, w_026_180, w_026_187, w_026_188, w_026_189, w_026_192, w_026_193, w_026_197, w_026_201, w_026_204, w_026_206, w_026_209, w_026_210, w_026_212, w_026_213, w_026_214, w_026_219, w_026_227, w_026_230, w_026_232, w_026_242, w_026_248, w_026_250, w_026_251, w_026_256, w_026_260, w_026_266, w_026_268, w_026_276, w_026_280, w_026_283, w_026_287, w_026_294, w_026_302, w_026_305, w_026_316, w_026_326, w_026_328, w_026_332, w_026_334, w_026_341, w_026_342, w_026_345, w_026_346, w_026_355, w_026_359, w_026_361, w_026_362, w_026_363, w_026_367, w_026_370, w_026_372, w_026_375, w_026_377, w_026_378, w_026_384, w_026_386, w_026_387, w_026_389, w_026_392;
  wire w_027_001, w_027_004, w_027_005, w_027_006, w_027_007, w_027_008, w_027_009, w_027_010, w_027_011, w_027_014, w_027_018, w_027_019, w_027_020, w_027_022, w_027_025, w_027_027, w_027_028, w_027_030, w_027_031, w_027_032, w_027_033, w_027_035, w_027_039, w_027_041, w_027_042, w_027_057, w_027_060, w_027_063, w_027_064, w_027_067, w_027_069, w_027_070, w_027_074, w_027_075, w_027_076, w_027_080, w_027_086, w_027_088, w_027_091, w_027_101, w_027_104, w_027_108, w_027_111, w_027_112, w_027_114, w_027_115, w_027_120, w_027_123, w_027_128, w_027_133, w_027_134, w_027_135, w_027_138, w_027_141, w_027_147, w_027_150, w_027_152, w_027_153, w_027_154, w_027_155, w_027_163, w_027_165, w_027_166, w_027_168, w_027_169, w_027_172, w_027_175, w_027_178, w_027_183, w_027_184, w_027_185, w_027_186, w_027_194, w_027_196, w_027_198, w_027_199, w_027_201, w_027_203, w_027_209, w_027_211, w_027_215, w_027_217, w_027_218, w_027_226, w_027_228, w_027_232, w_027_235, w_027_237, w_027_239, w_027_240, w_027_241, w_027_242, w_027_249, w_027_251, w_027_256, w_027_257, w_027_258, w_027_262, w_027_263, w_027_264, w_027_268, w_027_275, w_027_278, w_027_280, w_027_282, w_027_287, w_027_295, w_027_299, w_027_312, w_027_313, w_027_321, w_027_324, w_027_325, w_027_328, w_027_329, w_027_331, w_027_332, w_027_337, w_027_339, w_027_341, w_027_347, w_027_348, w_027_354, w_027_355, w_027_357, w_027_359, w_027_362, w_027_366, w_027_367, w_027_370, w_027_372, w_027_378, w_027_382, w_027_389, w_027_394, w_027_400, w_027_403, w_027_404, w_027_412, w_027_416, w_027_426, w_027_427, w_027_431, w_027_438, w_027_439, w_027_443, w_027_444, w_027_449, w_027_452;
  wire w_028_000, w_028_001, w_028_004, w_028_005, w_028_006, w_028_008, w_028_009, w_028_011, w_028_013, w_028_014, w_028_015, w_028_016, w_028_017, w_028_019, w_028_029, w_028_032, w_028_035, w_028_039, w_028_040, w_028_041, w_028_042, w_028_047, w_028_048, w_028_049, w_028_052, w_028_056, w_028_058, w_028_060, w_028_070, w_028_073, w_028_074, w_028_076, w_028_082, w_028_083, w_028_084, w_028_085, w_028_087, w_028_096, w_028_100, w_028_108, w_028_109, w_028_115, w_028_118, w_028_119, w_028_123, w_028_128, w_028_129, w_028_130, w_028_132, w_028_144, w_028_149, w_028_151, w_028_159, w_028_171, w_028_174, w_028_184, w_028_187, w_028_188, w_028_197, w_028_199, w_028_200, w_028_201, w_028_205, w_028_206, w_028_208, w_028_215, w_028_216, w_028_221, w_028_232, w_028_236, w_028_237, w_028_239, w_028_241, w_028_254, w_028_255, w_028_258, w_028_262, w_028_266, w_028_267, w_028_268, w_028_270, w_028_277, w_028_284, w_028_290, w_028_292, w_028_296, w_028_299, w_028_305, w_028_308, w_028_309, w_028_313, w_028_316, w_028_323, w_028_324, w_028_325, w_028_332, w_028_334, w_028_335, w_028_339, w_028_341, w_028_345, w_028_348, w_028_350, w_028_353, w_028_355, w_028_356, w_028_360, w_028_364, w_028_370, w_028_379, w_028_381, w_028_382, w_028_386, w_028_395, w_028_397;
  wire w_029_001, w_029_006, w_029_010, w_029_012, w_029_013, w_029_014, w_029_017, w_029_019, w_029_024, w_029_025, w_029_028, w_029_029, w_029_031, w_029_039, w_029_040, w_029_043, w_029_044, w_029_045, w_029_047, w_029_052, w_029_057, w_029_059, w_029_061, w_029_063, w_029_067, w_029_068, w_029_071, w_029_073, w_029_075, w_029_077, w_029_078, w_029_080, w_029_082, w_029_083, w_029_086, w_029_095, w_029_096, w_029_097, w_029_098, w_029_099, w_029_107, w_029_111, w_029_112, w_029_113, w_029_115, w_029_116, w_029_118, w_029_119, w_029_121, w_029_122, w_029_124, w_029_128, w_029_130, w_029_133, w_029_136, w_029_137, w_029_139, w_029_141, w_029_142, w_029_147, w_029_149, w_029_151, w_029_152, w_029_153, w_029_154, w_029_157, w_029_160, w_029_161, w_029_163, w_029_166, w_029_167, w_029_172, w_029_173, w_029_175, w_029_176, w_029_177, w_029_178, w_029_179, w_029_181, w_029_182, w_029_184, w_029_186, w_029_187, w_029_188, w_029_189, w_029_192, w_029_194, w_029_195, w_029_197, w_029_198, w_029_201, w_029_202, w_029_204, w_029_213, w_029_215, w_029_217, w_029_220, w_029_221, w_029_222, w_029_223, w_029_225, w_029_229, w_029_231, w_029_232, w_029_233, w_029_234, w_029_237, w_029_240, w_029_241, w_029_242, w_029_243, w_029_245, w_029_246, w_029_247, w_029_249, w_029_250, w_029_251, w_029_252, w_029_253, w_029_254, w_029_255, w_029_256, w_029_260, w_029_261, w_029_262, w_029_263, w_029_265;
  wire w_030_002, w_030_003, w_030_006, w_030_010, w_030_012, w_030_016, w_030_017, w_030_019, w_030_022, w_030_024, w_030_026, w_030_027, w_030_029, w_030_030, w_030_031, w_030_035, w_030_040, w_030_041, w_030_043, w_030_045, w_030_047, w_030_049, w_030_051, w_030_053, w_030_054, w_030_055, w_030_056, w_030_059, w_030_060, w_030_061, w_030_062, w_030_065, w_030_066, w_030_067, w_030_068, w_030_071, w_030_072, w_030_076, w_030_077, w_030_078, w_030_080, w_030_081, w_030_085, w_030_086, w_030_087, w_030_088, w_030_089, w_030_090, w_030_091, w_030_093, w_030_096, w_030_097, w_030_098, w_030_099, w_030_101, w_030_107, w_030_113, w_030_116, w_030_118, w_030_119, w_030_122, w_030_124, w_030_128, w_030_129, w_030_132, w_030_133, w_030_135, w_030_136, w_030_137, w_030_138, w_030_139, w_030_140, w_030_144, w_030_146, w_030_147, w_030_148, w_030_150, w_030_151, w_030_157, w_030_160, w_030_170, w_030_172, w_030_175, w_030_176, w_030_178, w_030_180, w_030_184, w_030_185, w_030_186, w_030_188, w_030_189, w_030_191, w_030_193, w_030_196, w_030_199;
  wire w_031_000, w_031_001, w_031_002, w_031_003, w_031_004, w_031_005, w_031_006, w_031_007, w_031_008, w_031_010, w_031_011, w_031_012, w_031_013, w_031_014, w_031_015, w_031_016, w_031_017, w_031_018, w_031_019, w_031_020, w_031_021, w_031_022, w_031_023, w_031_024, w_031_025, w_031_027, w_031_029, w_031_030, w_031_031, w_031_032, w_031_033, w_031_034, w_031_036, w_031_037, w_031_038, w_031_040, w_031_041, w_031_042, w_031_043, w_031_044, w_031_045, w_031_046, w_031_048, w_031_049, w_031_050, w_031_051, w_031_052, w_031_053, w_031_054, w_031_055, w_031_056, w_031_057, w_031_058, w_031_061, w_031_062, w_031_063, w_031_064, w_031_065, w_031_066, w_031_067;
  wire w_032_000, w_032_002, w_032_003, w_032_004, w_032_006, w_032_008, w_032_011, w_032_013, w_032_014, w_032_015, w_032_018, w_032_019, w_032_022, w_032_023, w_032_025, w_032_026, w_032_027, w_032_030, w_032_034, w_032_035, w_032_037, w_032_039, w_032_041, w_032_042, w_032_043, w_032_045, w_032_048, w_032_049, w_032_051, w_032_052, w_032_053, w_032_054, w_032_055, w_032_058, w_032_059, w_032_061, w_032_065, w_032_066, w_032_068, w_032_069, w_032_070, w_032_071, w_032_072, w_032_073, w_032_074, w_032_077, w_032_078, w_032_079, w_032_081, w_032_082, w_032_084, w_032_085, w_032_087, w_032_090, w_032_091, w_032_096, w_032_098, w_032_102, w_032_103, w_032_104, w_032_106, w_032_108, w_032_110, w_032_114, w_032_115, w_032_120, w_032_121, w_032_122, w_032_123, w_032_124, w_032_127, w_032_132, w_032_137, w_032_139, w_032_141, w_032_142, w_032_143, w_032_145, w_032_148, w_032_153, w_032_154, w_032_158, w_032_160, w_032_165, w_032_167, w_032_169, w_032_171, w_032_172, w_032_176, w_032_177, w_032_179, w_032_181, w_032_183, w_032_184, w_032_187, w_032_188, w_032_190, w_032_195;
  wire w_033_000, w_033_001, w_033_002, w_033_003, w_033_004, w_033_005, w_033_007, w_033_008, w_033_009, w_033_010, w_033_011, w_033_012, w_033_013, w_033_014, w_033_015, w_033_016, w_033_018, w_033_019, w_033_020, w_033_021, w_033_022, w_033_023, w_033_024, w_033_025, w_033_026, w_033_027, w_033_028, w_033_029, w_033_030, w_033_031, w_033_032, w_033_033, w_033_034, w_033_035, w_033_037, w_033_038, w_033_039, w_033_040, w_033_042, w_033_043, w_033_044, w_033_045, w_033_046, w_033_047, w_033_048, w_033_050, w_033_051, w_033_052, w_033_053, w_033_054, w_033_055, w_033_056, w_033_057, w_033_058;
  wire w_034_003, w_034_006, w_034_007, w_034_008, w_034_011, w_034_014, w_034_016, w_034_021, w_034_022, w_034_025, w_034_027, w_034_030, w_034_031, w_034_032, w_034_036, w_034_037, w_034_042, w_034_043, w_034_045, w_034_048, w_034_052, w_034_053, w_034_056, w_034_057, w_034_058, w_034_059, w_034_060, w_034_061, w_034_062, w_034_066, w_034_067, w_034_075, w_034_076, w_034_077, w_034_080, w_034_081, w_034_084, w_034_085, w_034_088, w_034_089, w_034_093, w_034_095, w_034_097, w_034_098, w_034_100, w_034_101, w_034_104, w_034_108, w_034_121, w_034_122, w_034_124, w_034_129, w_034_138, w_034_139, w_034_145, w_034_146, w_034_150, w_034_152, w_034_154, w_034_155, w_034_165, w_034_166, w_034_170, w_034_172, w_034_177, w_034_179, w_034_182, w_034_187, w_034_191, w_034_192, w_034_193, w_034_194, w_034_195, w_034_196, w_034_199, w_034_200, w_034_202, w_034_203, w_034_205, w_034_206, w_034_210, w_034_213, w_034_215, w_034_219, w_034_221, w_034_222, w_034_223, w_034_224, w_034_238, w_034_240, w_034_247, w_034_252, w_034_254, w_034_257, w_034_259, w_034_262, w_034_265, w_034_267, w_034_271, w_034_272, w_034_276, w_034_278, w_034_281;
  wire w_035_000, w_035_001, w_035_002, w_035_004, w_035_005, w_035_006, w_035_007, w_035_008, w_035_009, w_035_010, w_035_011, w_035_013, w_035_014, w_035_015, w_035_016, w_035_017, w_035_018, w_035_021, w_035_023, w_035_024, w_035_025, w_035_027, w_035_028, w_035_029, w_035_031, w_035_032, w_035_034, w_035_035, w_035_036, w_035_037, w_035_038, w_035_039, w_035_040, w_035_041, w_035_045, w_035_046, w_035_047, w_035_048, w_035_049, w_035_050, w_035_051, w_035_054, w_035_056, w_035_057, w_035_061, w_035_062, w_035_065, w_035_066, w_035_068, w_035_069, w_035_071, w_035_075, w_035_077, w_035_078, w_035_079, w_035_080, w_035_083, w_035_084, w_035_085, w_035_086, w_035_088, w_035_089, w_035_090, w_035_094, w_035_096, w_035_097, w_035_100, w_035_101, w_035_107, w_035_108, w_035_109;
  wire w_036_005, w_036_006, w_036_008, w_036_016, w_036_017, w_036_025, w_036_027, w_036_028, w_036_030, w_036_031, w_036_034, w_036_042, w_036_043, w_036_044, w_036_045, w_036_046, w_036_056, w_036_058, w_036_060, w_036_061, w_036_065, w_036_067, w_036_073, w_036_077, w_036_078, w_036_079, w_036_080, w_036_081, w_036_084, w_036_087, w_036_093, w_036_094, w_036_095, w_036_098, w_036_099, w_036_101, w_036_105, w_036_108, w_036_113, w_036_118, w_036_120, w_036_127, w_036_128, w_036_129, w_036_131, w_036_141, w_036_143, w_036_147, w_036_152, w_036_155, w_036_157, w_036_163, w_036_165, w_036_166, w_036_168, w_036_169, w_036_171, w_036_175, w_036_179, w_036_181, w_036_184, w_036_188, w_036_190, w_036_195, w_036_196, w_036_200, w_036_201, w_036_202, w_036_204, w_036_205, w_036_209, w_036_216, w_036_219, w_036_227, w_036_229, w_036_234, w_036_260, w_036_261, w_036_272, w_036_278;
  wire w_037_001, w_037_002, w_037_004, w_037_010, w_037_011, w_037_013, w_037_014, w_037_015, w_037_018, w_037_020, w_037_021, w_037_022, w_037_023, w_037_024, w_037_029, w_037_030, w_037_031, w_037_032, w_037_035, w_037_036, w_037_037, w_037_038, w_037_041, w_037_042, w_037_043, w_037_047, w_037_048, w_037_049, w_037_050, w_037_052, w_037_053, w_037_057, w_037_058, w_037_059, w_037_060, w_037_064, w_037_065, w_037_066, w_037_067, w_037_068, w_037_069, w_037_072, w_037_075, w_037_076, w_037_078, w_037_081, w_037_084, w_037_085, w_037_086, w_037_087, w_037_089, w_037_090, w_037_091, w_037_093, w_037_097, w_037_100, w_037_101, w_037_114, w_037_115, w_037_116, w_037_117, w_037_118, w_037_119, w_037_120, w_037_121, w_037_122, w_037_124, w_037_125, w_037_126, w_037_127, w_037_128, w_037_130, w_037_132, w_037_138, w_037_140, w_037_142, w_037_143, w_037_144, w_037_149;
  wire w_038_000, w_038_001, w_038_002, w_038_005, w_038_007, w_038_008, w_038_009, w_038_010, w_038_011, w_038_012, w_038_013, w_038_014, w_038_016, w_038_019, w_038_020, w_038_021, w_038_022, w_038_023, w_038_024, w_038_026, w_038_028, w_038_030, w_038_031, w_038_032, w_038_035, w_038_037, w_038_040, w_038_041, w_038_044, w_038_046, w_038_047, w_038_049, w_038_051, w_038_054, w_038_055, w_038_056, w_038_058, w_038_062, w_038_064, w_038_066, w_038_067, w_038_068, w_038_069, w_038_070, w_038_073, w_038_074, w_038_075, w_038_077, w_038_079, w_038_080, w_038_081, w_038_082, w_038_086, w_038_087, w_038_088, w_038_089, w_038_093, w_038_094, w_038_096, w_038_099;
  wire w_039_001, w_039_002, w_039_014, w_039_024, w_039_040, w_039_046, w_039_048, w_039_056, w_039_057, w_039_060, w_039_063, w_039_067, w_039_077, w_039_080, w_039_083, w_039_085, w_039_089, w_039_093, w_039_100, w_039_103, w_039_104, w_039_107, w_039_108, w_039_109, w_039_111, w_039_113, w_039_117, w_039_130, w_039_136, w_039_145, w_039_146, w_039_151, w_039_153, w_039_158, w_039_160, w_039_176, w_039_177, w_039_182, w_039_191, w_039_198, w_039_204, w_039_212, w_039_215, w_039_216, w_039_220, w_039_221, w_039_223, w_039_224, w_039_225, w_039_237, w_039_240, w_039_241, w_039_250, w_039_254, w_039_268, w_039_270, w_039_272, w_039_274, w_039_278, w_039_292, w_039_295, w_039_306, w_039_309, w_039_331, w_039_334, w_039_337, w_039_338, w_039_343, w_039_344, w_039_346, w_039_348, w_039_354, w_039_356, w_039_357, w_039_364, w_039_366, w_039_367, w_039_370, w_039_374, w_039_376, w_039_381, w_039_394, w_039_395, w_039_396, w_039_397, w_039_400, w_039_402, w_039_404, w_039_421, w_039_435, w_039_441, w_039_448, w_039_451, w_039_454, w_039_463, w_039_475, w_039_483, w_039_494, w_039_496, w_039_499, w_039_500, w_039_501, w_039_502, w_039_503, w_039_504, w_039_505, w_039_506, w_039_507, w_039_508, w_039_509, w_039_513, w_039_514, w_039_515, w_039_516, w_039_517, w_039_518, w_039_519, w_039_520, w_039_522;
  wire w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006;
  wire w_041_000, w_041_003, w_041_004, w_041_006, w_041_007, w_041_011, w_041_013, w_041_022, w_041_024, w_041_025, w_041_031, w_041_033, w_041_036, w_041_037, w_041_038, w_041_039, w_041_040, w_041_048, w_041_052, w_041_056, w_041_058, w_041_059, w_041_064, w_041_065, w_041_071, w_041_072, w_041_073, w_041_075, w_041_077, w_041_081, w_041_087, w_041_088, w_041_091, w_041_096, w_041_098, w_041_099, w_041_101, w_041_109, w_041_113, w_041_114, w_041_122, w_041_125, w_041_128, w_041_129, w_041_130, w_041_132, w_041_135, w_041_136, w_041_138, w_041_139, w_041_140, w_041_141, w_041_142, w_041_147, w_041_150, w_041_151, w_041_154, w_041_155, w_041_160, w_041_164, w_041_167, w_041_168, w_041_169, w_041_173, w_041_175, w_041_182, w_041_185, w_041_186, w_041_195, w_041_207, w_041_208, w_041_211, w_041_214, w_041_217, w_041_222, w_041_223, w_041_228, w_041_235, w_041_241, w_041_255, w_041_260, w_041_271, w_041_288, w_041_291, w_041_295, w_041_298, w_041_300;
  wire w_042_001, w_042_002, w_042_005, w_042_013, w_042_016, w_042_033, w_042_040, w_042_044, w_042_047, w_042_051, w_042_054, w_042_055, w_042_058, w_042_065, w_042_067, w_042_072, w_042_073, w_042_075, w_042_077, w_042_078, w_042_082, w_042_084, w_042_088, w_042_092, w_042_094, w_042_096, w_042_099, w_042_101, w_042_102, w_042_106, w_042_108, w_042_110, w_042_111, w_042_113, w_042_120, w_042_121, w_042_126, w_042_131, w_042_133, w_042_134, w_042_138, w_042_142, w_042_145, w_042_152, w_042_154, w_042_158, w_042_160, w_042_163, w_042_166, w_042_169, w_042_170, w_042_177, w_042_178, w_042_183, w_042_187, w_042_188, w_042_189, w_042_193, w_042_196, w_042_199, w_042_200, w_042_202, w_042_206, w_042_212, w_042_217, w_042_221, w_042_223, w_042_232, w_042_234, w_042_250, w_042_255, w_042_265, w_042_270, w_042_275;
  wire w_043_000, w_043_006, w_043_007, w_043_011, w_043_014, w_043_016, w_043_019, w_043_022, w_043_026, w_043_029, w_043_032, w_043_035, w_043_037, w_043_043, w_043_052, w_043_056, w_043_059, w_043_060, w_043_063, w_043_064, w_043_065, w_043_069, w_043_071, w_043_077, w_043_080, w_043_082, w_043_089, w_043_092, w_043_093, w_043_094, w_043_099, w_043_101, w_043_103, w_043_111, w_043_113, w_043_119, w_043_121, w_043_129, w_043_139, w_043_141, w_043_143, w_043_156, w_043_161, w_043_171, w_043_174, w_043_179, w_043_183, w_043_190, w_043_192, w_043_198, w_043_202, w_043_206, w_043_211, w_043_212, w_043_215, w_043_217, w_043_218, w_043_222, w_043_225, w_043_226, w_043_227, w_043_230, w_043_233, w_043_237, w_043_238, w_043_241, w_043_242;
  wire w_044_001, w_044_007, w_044_008, w_044_013, w_044_014, w_044_018, w_044_021, w_044_023, w_044_025, w_044_028, w_044_032, w_044_034, w_044_036, w_044_037, w_044_038, w_044_048, w_044_049, w_044_050, w_044_053, w_044_055, w_044_059, w_044_062, w_044_070, w_044_073, w_044_074, w_044_075, w_044_087, w_044_091, w_044_094, w_044_101, w_044_108, w_044_109, w_044_110, w_044_112, w_044_119, w_044_120, w_044_127, w_044_130, w_044_133, w_044_136, w_044_140, w_044_146, w_044_151, w_044_153, w_044_154, w_044_157, w_044_158, w_044_161, w_044_163, w_044_169, w_044_171, w_044_172, w_044_184, w_044_193, w_044_210, w_044_212, w_044_216, w_044_220, w_044_227, w_044_237, w_044_240, w_044_242, w_044_245, w_044_258, w_044_259, w_044_264, w_044_269, w_044_275, w_044_277, w_044_281, w_044_282, w_044_295, w_044_297, w_044_301, w_044_302, w_044_307, w_044_323, w_044_326;
  wire w_045_001, w_045_004, w_045_005, w_045_008, w_045_009, w_045_010, w_045_015, w_045_018, w_045_026, w_045_036, w_045_038, w_045_039, w_045_065, w_045_066, w_045_069, w_045_082, w_045_090, w_045_092, w_045_094, w_045_096, w_045_099, w_045_103, w_045_104, w_045_106, w_045_112, w_045_114, w_045_115, w_045_118, w_045_119, w_045_125, w_045_132, w_045_135, w_045_136, w_045_137, w_045_139, w_045_150, w_045_152, w_045_170, w_045_171, w_045_174, w_045_177, w_045_180, w_045_182, w_045_183, w_045_184, w_045_185, w_045_193, w_045_199, w_045_201, w_045_210, w_045_216, w_045_229, w_045_231, w_045_241, w_045_250, w_045_257, w_045_276, w_045_283, w_045_284;
  wire w_046_004, w_046_005, w_046_006, w_046_007, w_046_008, w_046_010, w_046_011, w_046_015, w_046_016, w_046_021, w_046_023, w_046_024, w_046_026, w_046_027, w_046_028, w_046_031, w_046_032, w_046_035, w_046_037, w_046_039, w_046_040, w_046_043, w_046_044, w_046_045, w_046_047, w_046_048, w_046_053, w_046_056, w_046_060, w_046_061, w_046_062, w_046_063, w_046_067, w_046_084, w_046_086, w_046_090, w_046_094, w_046_097, w_046_107, w_046_108, w_046_113, w_046_114, w_046_115, w_046_118, w_046_119, w_046_122, w_046_125, w_046_126, w_046_127, w_046_132, w_046_134, w_046_138, w_046_145, w_046_148, w_046_150, w_046_151, w_046_161, w_046_165, w_046_166, w_046_170, w_046_171, w_046_173, w_046_174, w_046_178, w_046_179, w_046_180, w_046_182, w_046_183, w_046_185, w_046_192, w_046_198, w_046_208, w_046_210, w_046_211, w_046_216, w_046_218, w_046_221;
  wire w_047_001, w_047_007, w_047_013, w_047_015, w_047_022, w_047_023, w_047_030, w_047_032, w_047_036, w_047_038, w_047_044, w_047_045, w_047_046, w_047_050, w_047_053, w_047_054, w_047_062, w_047_064, w_047_089, w_047_090, w_047_102, w_047_103, w_047_113, w_047_134, w_047_137, w_047_141, w_047_151, w_047_152, w_047_154, w_047_162, w_047_164, w_047_165, w_047_173, w_047_174, w_047_175, w_047_179, w_047_183, w_047_185, w_047_196, w_047_201, w_047_202, w_047_207, w_047_216, w_047_224, w_047_228, w_047_229, w_047_230, w_047_231, w_047_233, w_047_234, w_047_235, w_047_251, w_047_253, w_047_256, w_047_258, w_047_259, w_047_267, w_047_274, w_047_276, w_047_278, w_047_279, w_047_286, w_047_288, w_047_291, w_047_292, w_047_293, w_047_306, w_047_310, w_047_316, w_047_317, w_047_318, w_047_322, w_047_329, w_047_330, w_047_336, w_047_339, w_047_341, w_047_350, w_047_354, w_047_367, w_047_368, w_047_390, w_047_397, w_047_400, w_047_405, w_047_415, w_047_416, w_047_422;
  wire w_048_000, w_048_001, w_048_003, w_048_012, w_048_014, w_048_019, w_048_020, w_048_021, w_048_022, w_048_026, w_048_029, w_048_033, w_048_050, w_048_054, w_048_055, w_048_056, w_048_061, w_048_064, w_048_071, w_048_072, w_048_074, w_048_079, w_048_081, w_048_083, w_048_085, w_048_087, w_048_097, w_048_100, w_048_103, w_048_104, w_048_107, w_048_109, w_048_117, w_048_118, w_048_119, w_048_128, w_048_132, w_048_133, w_048_137, w_048_143, w_048_147, w_048_149, w_048_169, w_048_171, w_048_184, w_048_187, w_048_190, w_048_193, w_048_196, w_048_207, w_048_209, w_048_211, w_048_216, w_048_233, w_048_234, w_048_247, w_048_255, w_048_265, w_048_268, w_048_271, w_048_279, w_048_280, w_048_281, w_048_284, w_048_285, w_048_303, w_048_304, w_048_314, w_048_317, w_048_342, w_048_347, w_048_355, w_048_366;
  wire w_049_000, w_049_002, w_049_003, w_049_008, w_049_012, w_049_023, w_049_025, w_049_030, w_049_038, w_049_044, w_049_047, w_049_060, w_049_065, w_049_066, w_049_070, w_049_071, w_049_074, w_049_076, w_049_079, w_049_087, w_049_090, w_049_091, w_049_100, w_049_107, w_049_108, w_049_113, w_049_121, w_049_137, w_049_139, w_049_149, w_049_165, w_049_166, w_049_173, w_049_174, w_049_179, w_049_182, w_049_185, w_049_189, w_049_191, w_049_200, w_049_201, w_049_218, w_049_219, w_049_231, w_049_244, w_049_250, w_049_262, w_049_266, w_049_272, w_049_273, w_049_277, w_049_285, w_049_297, w_049_301, w_049_307, w_049_320, w_049_323, w_049_329, w_049_333, w_049_338, w_049_343, w_049_347, w_049_361, w_049_377, w_049_380, w_049_383, w_049_388, w_049_400, w_049_401, w_049_403;
  wire w_050_001, w_050_002, w_050_003, w_050_007, w_050_008, w_050_009, w_050_010, w_050_014, w_050_015, w_050_016, w_050_017, w_050_022, w_050_026, w_050_030, w_050_034, w_050_035, w_050_038, w_050_039, w_050_042, w_050_043, w_050_045, w_050_046, w_050_047, w_050_051, w_050_052, w_050_054, w_050_055, w_050_057, w_050_058, w_050_060, w_050_063, w_050_067, w_050_070, w_050_073, w_050_087, w_050_096, w_050_102, w_050_106, w_050_111, w_050_112, w_050_113, w_050_117, w_050_121, w_050_124, w_050_125, w_050_126, w_050_128, w_050_136, w_050_138, w_050_142, w_050_146, w_050_149, w_050_152, w_050_155, w_050_161, w_050_172, w_050_173, w_050_174, w_050_175, w_050_176, w_050_180, w_050_182, w_050_184, w_050_187, w_050_188, w_050_192, w_050_193, w_050_198, w_050_199, w_050_204;
  wire w_051_001, w_051_002, w_051_003, w_051_008, w_051_010, w_051_016, w_051_017, w_051_018, w_051_023, w_051_026, w_051_028, w_051_031, w_051_033, w_051_035, w_051_041, w_051_042, w_051_045, w_051_046, w_051_056, w_051_060, w_051_076, w_051_078, w_051_081, w_051_085, w_051_094, w_051_095, w_051_097, w_051_098, w_051_101, w_051_104, w_051_107, w_051_110, w_051_117, w_051_119, w_051_124, w_051_128, w_051_130, w_051_132, w_051_146, w_051_151, w_051_153, w_051_154, w_051_159, w_051_164, w_051_165, w_051_172, w_051_181, w_051_182, w_051_197, w_051_198, w_051_210, w_051_211, w_051_218, w_051_221, w_051_223, w_051_226, w_051_238, w_051_246, w_051_253, w_051_260, w_051_266, w_051_286, w_051_306, w_051_313;
  wire w_052_004, w_052_005, w_052_006, w_052_007, w_052_008, w_052_009, w_052_012, w_052_013, w_052_015, w_052_016, w_052_017, w_052_018, w_052_019, w_052_020, w_052_022, w_052_023, w_052_027, w_052_033, w_052_034, w_052_035, w_052_036, w_052_038, w_052_039, w_052_040, w_052_047, w_052_048, w_052_049, w_052_051, w_052_054, w_052_056, w_052_058, w_052_061, w_052_066, w_052_068, w_052_071, w_052_084, w_052_085, w_052_086, w_052_095, w_052_097, w_052_098, w_052_101, w_052_103, w_052_104, w_052_110, w_052_112, w_052_113, w_052_115, w_052_116;
  wire w_053_000, w_053_001, w_053_002, w_053_003, w_053_004, w_053_005, w_053_006, w_053_007, w_053_009, w_053_011, w_053_013, w_053_014, w_053_015, w_053_016, w_053_018, w_053_019, w_053_021, w_053_022, w_053_023, w_053_025, w_053_026, w_053_027, w_053_028, w_053_029, w_053_031, w_053_033, w_053_034, w_053_035, w_053_037, w_053_039;
  wire w_054_000, w_054_003, w_054_005, w_054_012, w_054_013, w_054_014, w_054_015, w_054_018, w_054_020, w_054_023, w_054_029, w_054_030, w_054_031, w_054_034, w_054_038, w_054_040, w_054_042, w_054_043, w_054_044, w_054_048, w_054_051, w_054_054, w_054_055, w_054_056, w_054_057, w_054_063, w_054_064, w_054_068, w_054_070, w_054_073, w_054_074, w_054_081, w_054_083, w_054_084, w_054_088, w_054_089, w_054_090, w_054_097, w_054_100, w_054_101, w_054_106, w_054_110, w_054_113, w_054_115, w_054_118, w_054_125, w_054_134, w_054_137, w_054_146, w_054_165, w_054_166, w_054_170, w_054_172, w_054_177, w_054_178, w_054_191, w_054_199, w_054_204, w_054_205, w_054_208, w_054_210, w_054_211;
  wire w_055_000, w_055_001, w_055_002, w_055_005, w_055_011, w_055_012, w_055_016, w_055_018, w_055_019, w_055_022, w_055_028, w_055_029, w_055_031, w_055_033, w_055_035, w_055_036, w_055_037, w_055_039, w_055_040, w_055_043, w_055_045, w_055_046, w_055_047, w_055_048, w_055_049, w_055_051, w_055_052, w_055_053, w_055_055, w_055_056, w_055_059, w_055_064, w_055_065, w_055_068, w_055_069, w_055_071, w_055_072, w_055_074, w_055_075, w_055_076, w_055_077, w_055_078, w_055_079, w_055_083, w_055_085, w_055_086;
  wire w_056_003, w_056_008, w_056_010, w_056_015, w_056_020, w_056_026, w_056_036, w_056_043, w_056_046, w_056_047, w_056_048, w_056_050, w_056_053, w_056_054, w_056_056, w_056_058, w_056_063, w_056_068, w_056_071, w_056_074, w_056_076, w_056_078, w_056_087, w_056_092, w_056_093, w_056_100, w_056_102, w_056_105, w_056_106, w_056_109, w_056_110, w_056_111, w_056_118, w_056_121, w_056_122, w_056_131, w_056_137, w_056_138, w_056_139, w_056_141, w_056_142, w_056_143, w_056_146, w_056_147, w_056_148, w_056_149, w_056_151, w_056_162, w_056_163, w_056_164, w_056_169, w_056_170, w_056_175, w_056_176, w_056_177;
  wire w_057_001, w_057_002, w_057_003, w_057_004, w_057_005, w_057_006, w_057_007, w_057_008, w_057_010, w_057_011, w_057_012, w_057_015, w_057_016, w_057_018, w_057_019, w_057_020, w_057_021, w_057_022, w_057_023, w_057_024, w_057_027, w_057_028, w_057_030, w_057_031, w_057_033, w_057_034, w_057_035, w_057_036, w_057_037, w_057_039, w_057_041, w_057_044, w_057_046, w_057_048, w_057_049, w_057_050, w_057_051, w_057_052, w_057_053, w_057_054, w_057_056, w_057_057, w_057_058, w_057_059, w_057_060;
  wire w_058_000, w_058_001, w_058_005, w_058_007, w_058_010, w_058_012, w_058_014, w_058_016, w_058_017, w_058_020, w_058_021, w_058_023, w_058_024, w_058_025, w_058_027, w_058_031, w_058_032, w_058_034, w_058_035, w_058_037, w_058_038, w_058_040, w_058_041, w_058_047, w_058_048, w_058_051, w_058_052, w_058_056, w_058_058, w_058_059, w_058_062, w_058_068, w_058_072, w_058_073, w_058_074, w_058_075, w_058_076, w_058_079, w_058_081, w_058_083, w_058_084, w_058_086;
  wire w_059_004, w_059_018, w_059_025, w_059_028, w_059_032, w_059_041, w_059_046, w_059_056, w_059_063, w_059_072, w_059_077, w_059_095, w_059_100, w_059_120, w_059_121, w_059_133, w_059_148, w_059_158, w_059_159, w_059_168, w_059_169, w_059_191, w_059_195, w_059_199, w_059_211, w_059_216, w_059_217, w_059_223, w_059_233, w_059_237, w_059_255, w_059_256, w_059_260, w_059_262, w_059_264, w_059_267, w_059_269, w_059_272, w_059_280, w_059_284, w_059_288, w_059_293, w_059_297, w_059_317, w_059_318, w_059_322, w_059_337, w_059_341, w_059_344, w_059_346, w_059_348, w_059_351, w_059_358, w_059_359, w_059_390, w_059_403, w_059_415, w_059_438, w_059_440, w_059_444, w_059_445, w_059_461, w_059_478, w_059_484;
  wire w_060_009, w_060_010, w_060_011, w_060_017, w_060_020, w_060_023, w_060_027, w_060_032, w_060_033, w_060_040, w_060_045, w_060_047, w_060_049, w_060_050, w_060_055, w_060_060, w_060_064, w_060_065, w_060_089, w_060_096, w_060_111, w_060_117, w_060_124, w_060_125, w_060_135, w_060_142, w_060_144, w_060_153, w_060_166, w_060_174, w_060_179, w_060_184, w_060_187, w_060_194, w_060_220, w_060_226, w_060_242, w_060_260, w_060_267, w_060_268, w_060_290, w_060_295, w_060_303, w_060_315, w_060_322, w_060_334, w_060_344, w_060_370, w_060_379, w_060_432;
  wire w_061_000, w_061_008, w_061_014, w_061_023, w_061_024, w_061_025, w_061_027, w_061_032, w_061_039, w_061_041, w_061_047, w_061_050, w_061_062, w_061_066, w_061_072, w_061_094, w_061_114, w_061_117, w_061_126, w_061_127, w_061_130, w_061_144, w_061_160, w_061_170, w_061_174, w_061_178, w_061_190, w_061_199, w_061_207, w_061_208, w_061_212, w_061_213, w_061_222, w_061_224, w_061_236, w_061_242, w_061_247, w_061_249, w_061_265, w_061_268, w_061_271, w_061_275, w_061_284, w_061_297, w_061_304, w_061_309, w_061_314, w_061_330, w_061_334, w_061_337, w_061_356, w_061_367, w_061_373, w_061_376, w_061_383, w_061_391, w_061_405, w_061_406, w_061_412, w_061_421;
  wire w_062_000, w_062_002, w_062_003, w_062_004, w_062_005, w_062_006, w_062_007, w_062_008, w_062_009, w_062_010, w_062_011, w_062_012, w_062_013, w_062_015, w_062_016, w_062_018, w_062_019, w_062_020;
  wire w_063_003, w_063_005, w_063_006, w_063_010, w_063_011, w_063_013, w_063_020, w_063_022, w_063_024, w_063_025, w_063_026, w_063_028, w_063_030, w_063_036, w_063_043, w_063_047, w_063_056, w_063_057, w_063_062, w_063_074, w_063_076, w_063_078, w_063_079, w_063_089, w_063_091, w_063_097, w_063_106, w_063_111, w_063_113, w_063_114, w_063_117, w_063_118, w_063_122, w_063_123, w_063_139, w_063_141, w_063_150, w_063_159, w_063_165, w_063_171, w_063_174, w_063_179, w_063_197, w_063_200, w_063_206, w_063_208, w_063_218, w_063_222, w_063_223, w_063_226, w_063_228, w_063_232, w_063_256;
  wire w_064_000, w_064_001, w_064_002, w_064_003, w_064_006, w_064_007, w_064_009, w_064_011, w_064_014, w_064_015, w_064_017, w_064_018, w_064_020, w_064_022, w_064_023, w_064_024, w_064_030, w_064_031, w_064_032, w_064_034, w_064_035, w_064_039, w_064_044, w_064_045, w_064_046, w_064_047, w_064_052, w_064_053, w_064_058, w_064_060, w_064_070;
  wire w_065_007, w_065_009, w_065_010, w_065_014, w_065_019, w_065_021, w_065_024, w_065_027, w_065_029, w_065_032, w_065_035, w_065_036, w_065_039, w_065_041, w_065_042, w_065_050, w_065_055, w_065_057, w_065_070, w_065_072, w_065_079, w_065_084, w_065_093, w_065_094, w_065_104, w_065_105, w_065_109, w_065_110, w_065_112, w_065_121, w_065_124, w_065_126, w_065_133, w_065_136, w_065_151, w_065_158, w_065_159, w_065_182, w_065_185, w_065_191, w_065_202, w_065_210, w_065_214, w_065_219;
  wire w_066_002, w_066_003, w_066_006, w_066_013, w_066_014, w_066_031, w_066_036, w_066_038, w_066_060, w_066_067, w_066_072, w_066_074, w_066_080, w_066_097, w_066_098, w_066_108, w_066_111, w_066_113, w_066_116, w_066_117, w_066_126, w_066_128, w_066_131, w_066_135, w_066_145, w_066_150, w_066_154, w_066_160, w_066_163, w_066_168, w_066_169;
  wire w_067_000, w_067_001, w_067_003, w_067_004, w_067_006, w_067_007, w_067_008, w_067_009, w_067_014, w_067_015, w_067_016, w_067_017, w_067_020, w_067_022, w_067_023, w_067_025, w_067_026, w_067_029, w_067_030, w_067_031, w_067_032, w_067_033, w_067_035, w_067_036, w_067_039, w_067_040, w_067_044, w_067_045, w_067_050, w_067_051, w_067_055, w_067_056, w_067_059, w_067_060, w_067_061, w_067_062;
  wire w_068_000, w_068_002, w_068_003, w_068_006, w_068_009, w_068_011, w_068_012, w_068_014, w_068_016, w_068_020, w_068_022, w_068_025, w_068_032, w_068_036, w_068_040, w_068_042, w_068_046, w_068_048, w_068_051, w_068_053, w_068_055, w_068_058, w_068_066, w_068_070, w_068_076, w_068_080, w_068_087, w_068_090, w_068_093, w_068_097, w_068_099, w_068_100, w_068_103, w_068_119, w_068_129, w_068_136, w_068_138, w_068_139, w_068_146, w_068_149, w_068_150, w_068_151, w_068_155, w_068_156;
  wire w_069_000, w_069_006, w_069_008, w_069_009, w_069_012, w_069_015, w_069_017, w_069_023, w_069_026, w_069_028, w_069_031, w_069_037, w_069_040, w_069_054, w_069_058, w_069_063, w_069_064, w_069_065, w_069_068, w_069_069, w_069_085, w_069_089, w_069_091, w_069_097, w_069_106, w_069_108, w_069_109, w_069_112, w_069_125, w_069_128, w_069_130, w_069_132, w_069_134, w_069_144, w_069_147, w_069_149, w_069_157, w_069_158, w_069_160, w_069_165;
  wire w_070_000, w_070_002, w_070_003, w_070_004, w_070_005, w_070_007, w_070_009, w_070_017, w_070_018, w_070_022, w_070_024, w_070_031, w_070_032, w_070_034, w_070_040, w_070_041, w_070_042, w_070_046, w_070_047, w_070_048, w_070_053, w_070_055, w_070_058, w_070_059, w_070_061, w_070_065, w_070_067, w_070_068, w_070_070, w_070_072, w_070_074, w_070_076, w_070_079, w_070_081, w_070_084, w_070_085, w_070_087, w_070_090, w_070_091, w_070_094, w_070_095, w_070_099;
  wire w_071_004, w_071_005, w_071_010, w_071_020, w_071_036, w_071_046, w_071_055, w_071_088, w_071_089, w_071_094, w_071_104, w_071_116, w_071_122, w_071_147, w_071_148, w_071_156, w_071_158, w_071_169, w_071_185, w_071_191, w_071_193, w_071_205, w_071_211, w_071_212, w_071_214, w_071_225, w_071_235, w_071_270, w_071_289, w_071_294, w_071_295, w_071_299, w_071_311, w_071_321, w_071_347, w_071_348, w_071_352, w_071_354, w_071_358, w_071_362, w_071_367, w_071_389, w_071_394, w_071_395, w_071_410;
  wire w_072_006, w_072_007, w_072_008, w_072_011, w_072_014, w_072_018, w_072_020, w_072_022, w_072_031, w_072_034, w_072_042, w_072_045, w_072_048, w_072_050, w_072_053, w_072_054, w_072_058, w_072_064, w_072_065, w_072_067, w_072_068, w_072_073, w_072_074, w_072_075, w_072_080, w_072_084, w_072_086, w_072_088, w_072_096, w_072_097, w_072_100, w_072_102, w_072_104;
  wire w_073_001, w_073_007, w_073_009, w_073_010, w_073_012, w_073_014, w_073_016, w_073_017, w_073_021, w_073_023, w_073_026, w_073_027, w_073_028, w_073_036, w_073_039, w_073_040, w_073_041, w_073_043, w_073_044, w_073_046, w_073_069, w_073_072, w_073_074, w_073_078, w_073_099, w_073_101, w_073_111, w_073_117, w_073_123, w_073_125, w_073_129, w_073_132, w_073_133, w_073_138, w_073_149, w_073_172, w_073_173, w_073_176, w_073_181, w_073_187, w_073_189, w_073_191, w_073_218, w_073_222;
  wire w_074_000, w_074_001, w_074_002, w_074_003, w_074_004, w_074_005;
  wire w_075_018, w_075_020, w_075_021, w_075_022, w_075_024, w_075_025, w_075_038, w_075_040, w_075_041, w_075_042, w_075_047, w_075_053, w_075_054, w_075_056, w_075_067, w_075_070, w_075_074, w_075_080, w_075_081, w_075_084, w_075_087, w_075_089, w_075_091, w_075_093, w_075_094, w_075_095, w_075_099, w_075_100, w_075_103, w_075_109, w_075_113, w_075_118, w_075_121, w_075_122, w_075_124, w_075_130;
  wire w_076_000, w_076_008, w_076_009, w_076_011, w_076_013, w_076_018, w_076_020, w_076_021, w_076_023, w_076_026, w_076_029, w_076_031, w_076_033, w_076_039, w_076_042, w_076_045, w_076_056, w_076_058, w_076_060, w_076_062, w_076_065, w_076_068, w_076_069, w_076_070, w_076_075, w_076_077, w_076_078, w_076_085, w_076_086, w_076_093, w_076_094, w_076_095, w_076_097, w_076_102, w_076_104, w_076_107, w_076_115;
  wire w_077_012, w_077_024, w_077_029, w_077_037, w_077_038, w_077_052, w_077_053, w_077_057, w_077_061, w_077_083, w_077_085, w_077_086, w_077_099, w_077_101, w_077_104, w_077_109, w_077_113, w_077_117, w_077_120, w_077_123, w_077_125, w_077_135, w_077_142, w_077_148, w_077_153, w_077_156, w_077_157, w_077_162, w_077_164, w_077_174, w_077_184, w_077_185, w_077_191, w_077_201, w_077_236, w_077_246;
  wire w_078_000, w_078_001, w_078_002, w_078_006, w_078_011, w_078_012, w_078_013, w_078_019, w_078_028, w_078_032, w_078_041, w_078_050, w_078_053, w_078_055, w_078_057, w_078_062, w_078_063, w_078_066, w_078_067, w_078_071, w_078_074, w_078_078, w_078_081, w_078_086, w_078_090, w_078_091, w_078_094, w_078_099, w_078_104, w_078_107, w_078_116, w_078_117, w_078_123, w_078_126, w_078_136, w_078_142, w_078_143, w_078_144, w_078_160, w_078_161, w_078_163, w_078_164;
  wire w_079_007, w_079_013, w_079_020, w_079_021, w_079_028, w_079_040, w_079_047, w_079_065, w_079_133, w_079_141, w_079_158, w_079_170, w_079_181, w_079_193, w_079_197, w_079_199, w_079_219, w_079_224, w_079_235, w_079_237, w_079_247, w_079_256, w_079_257, w_079_267, w_079_304, w_079_320, w_079_328, w_079_342, w_079_362, w_079_401, w_079_402, w_079_407, w_079_422, w_079_432, w_079_434, w_079_452, w_079_453;
  wire w_080_000, w_080_001, w_080_003, w_080_004, w_080_005, w_080_007, w_080_009, w_080_011, w_080_012, w_080_013, w_080_014, w_080_015, w_080_016, w_080_017, w_080_018, w_080_019, w_080_020, w_080_021, w_080_023, w_080_024, w_080_025, w_080_028, w_080_031, w_080_032, w_080_035;
  wire w_081_001, w_081_003, w_081_004, w_081_008, w_081_010, w_081_011, w_081_012, w_081_017, w_081_018, w_081_020, w_081_025, w_081_026, w_081_027, w_081_029, w_081_030, w_081_034, w_081_035, w_081_037, w_081_038, w_081_039, w_081_044, w_081_053, w_081_058, w_081_061, w_081_064, w_081_069, w_081_073, w_081_074, w_081_082, w_081_083, w_081_084, w_081_087, w_081_088, w_081_089, w_081_090;
  wire w_082_000, w_082_002, w_082_005, w_082_007, w_082_015, w_082_018, w_082_027, w_082_032, w_082_038, w_082_039, w_082_053, w_082_059, w_082_088, w_082_101, w_082_103, w_082_106, w_082_113, w_082_122, w_082_125, w_082_126, w_082_134, w_082_141, w_082_144, w_082_158, w_082_188, w_082_196, w_082_197, w_082_212, w_082_221, w_082_234, w_082_242, w_082_270, w_082_275, w_082_316, w_082_338, w_082_340, w_082_341, w_082_342, w_082_343, w_082_344, w_082_345;
  wire w_083_000, w_083_002, w_083_003, w_083_004, w_083_011, w_083_012, w_083_013, w_083_022, w_083_023, w_083_025, w_083_031, w_083_035, w_083_046, w_083_056, w_083_061, w_083_079, w_083_083, w_083_084, w_083_090, w_083_098, w_083_103, w_083_105, w_083_107, w_083_108, w_083_111, w_083_119, w_083_123, w_083_125, w_083_159, w_083_160, w_083_171, w_083_177, w_083_179, w_083_188, w_083_195, w_083_205, w_083_208, w_083_212;
  wire w_084_000, w_084_005, w_084_006, w_084_010, w_084_012, w_084_020, w_084_026, w_084_030, w_084_031, w_084_037, w_084_051, w_084_053, w_084_055, w_084_062, w_084_076, w_084_085, w_084_086, w_084_103, w_084_111, w_084_113, w_084_114, w_084_122, w_084_132, w_084_136, w_084_137, w_084_163, w_084_176, w_084_201, w_084_207, w_084_214, w_084_237, w_084_261, w_084_268, w_084_270, w_084_286, w_084_288, w_084_321, w_084_327, w_084_337, w_084_342;
  wire w_085_002, w_085_017, w_085_021, w_085_027, w_085_036, w_085_044, w_085_055, w_085_057, w_085_060, w_085_065, w_085_066, w_085_079, w_085_098, w_085_108, w_085_113, w_085_119, w_085_124, w_085_127, w_085_138, w_085_139, w_085_144, w_085_158, w_085_159, w_085_177, w_085_182, w_085_197, w_085_206, w_085_223, w_085_236, w_085_244, w_085_246;
  wire w_086_001, w_086_007, w_086_010, w_086_024, w_086_026, w_086_038, w_086_042, w_086_043, w_086_047, w_086_052, w_086_055, w_086_068, w_086_070, w_086_073, w_086_084, w_086_092, w_086_095, w_086_100, w_086_102, w_086_103, w_086_107, w_086_120, w_086_123, w_086_133, w_086_140, w_086_148, w_086_149, w_086_157, w_086_158, w_086_160, w_086_161, w_086_165, w_086_188, w_086_192, w_086_195;
  wire w_087_004, w_087_019, w_087_027, w_087_038, w_087_039, w_087_061, w_087_062, w_087_067, w_087_074, w_087_082, w_087_083, w_087_104, w_087_130, w_087_138, w_087_142, w_087_147, w_087_148, w_087_149, w_087_178, w_087_188, w_087_217, w_087_218, w_087_240, w_087_279, w_087_281, w_087_314, w_087_322;
  wire w_088_012, w_088_021, w_088_030, w_088_031, w_088_041, w_088_061, w_088_107, w_088_119, w_088_123, w_088_132, w_088_136, w_088_163, w_088_199, w_088_245, w_088_252, w_088_270, w_088_278, w_088_315, w_088_335, w_088_336, w_088_392, w_088_397, w_088_409, w_088_410, w_088_421, w_088_435, w_088_445, w_088_454, w_088_455, w_088_456, w_088_460, w_088_461, w_088_462, w_088_463, w_088_464, w_088_465, w_088_466, w_088_467, w_088_468, w_088_469, w_088_471;
  wire w_089_001, w_089_007, w_089_026, w_089_031, w_089_032, w_089_035, w_089_046, w_089_074, w_089_090, w_089_092, w_089_096, w_089_101, w_089_103, w_089_120, w_089_138, w_089_180, w_089_189, w_089_193, w_089_217, w_089_221, w_089_243, w_089_264, w_089_273, w_089_288, w_089_305, w_089_307, w_089_380, w_089_400, w_089_404, w_089_416, w_089_429, w_089_431, w_089_442;
  wire w_090_012, w_090_017, w_090_019, w_090_064, w_090_068, w_090_076, w_090_079, w_090_087, w_090_089, w_090_101, w_090_111, w_090_120, w_090_128, w_090_139, w_090_141, w_090_163, w_090_177, w_090_186, w_090_190, w_090_194, w_090_215, w_090_221, w_090_228, w_090_249, w_090_256, w_090_262, w_090_281, w_090_283, w_090_287, w_090_288, w_090_290, w_090_298, w_090_301, w_090_317, w_090_319, w_090_326;
  wire w_091_003, w_091_040, w_091_045, w_091_052, w_091_054, w_091_070, w_091_076, w_091_077, w_091_109, w_091_123, w_091_124, w_091_135, w_091_152, w_091_168, w_091_174, w_091_189, w_091_225, w_091_235, w_091_243, w_091_253, w_091_254, w_091_258, w_091_260, w_091_264, w_091_289, w_091_326, w_091_342, w_091_354, w_091_371, w_091_411, w_091_417;
  wire w_092_005, w_092_009, w_092_014, w_092_016, w_092_017, w_092_023, w_092_026, w_092_032, w_092_033, w_092_035, w_092_038, w_092_045, w_092_049, w_092_064, w_092_065, w_092_068, w_092_073, w_092_074, w_092_076, w_092_085, w_092_087, w_092_094, w_092_107, w_092_109, w_092_112, w_092_123, w_092_129, w_092_156, w_092_166, w_092_171, w_092_176;
  wire w_093_000, w_093_004, w_093_009, w_093_018, w_093_024, w_093_034, w_093_039, w_093_053, w_093_064, w_093_072, w_093_095, w_093_101, w_093_107, w_093_110, w_093_111, w_093_115, w_093_143, w_093_152, w_093_161, w_093_186, w_093_208, w_093_209, w_093_216, w_093_246, w_093_258, w_093_264, w_093_266, w_093_269, w_093_272, w_093_276, w_093_281, w_093_293, w_093_295, w_093_318, w_093_329, w_093_346, w_093_348, w_093_351, w_093_364, w_093_365, w_093_371, w_093_378, w_093_426, w_093_427, w_093_428, w_093_429, w_093_430, w_093_434, w_093_435, w_093_436, w_093_437, w_093_438, w_093_439, w_093_440, w_093_441, w_093_442, w_093_443, w_093_444, w_093_445, w_093_447;
  wire w_094_003, w_094_010, w_094_014, w_094_023, w_094_028, w_094_033, w_094_045, w_094_049, w_094_062, w_094_081, w_094_147, w_094_155, w_094_166, w_094_171, w_094_199, w_094_229, w_094_319, w_094_320, w_094_357, w_094_393, w_094_416;
  wire w_095_000, w_095_001, w_095_002, w_095_010, w_095_014, w_095_016, w_095_017, w_095_023, w_095_026, w_095_030, w_095_036, w_095_037, w_095_038, w_095_044, w_095_048, w_095_049, w_095_051, w_095_052, w_095_058, w_095_061, w_095_064, w_095_066, w_095_067, w_095_073, w_095_080, w_095_084, w_095_089, w_095_091, w_095_094, w_095_099;
  wire w_096_004, w_096_009, w_096_010, w_096_017, w_096_018, w_096_020, w_096_022, w_096_024, w_096_026, w_096_027, w_096_030, w_096_033, w_096_038, w_096_039, w_096_046, w_096_054, w_096_059, w_096_086, w_096_095, w_096_102, w_096_106, w_096_127, w_096_134, w_096_136, w_096_145, w_096_146, w_096_147, w_096_150, w_096_151, w_096_154, w_096_155, w_096_165, w_096_174, w_096_176, w_096_184, w_096_197, w_096_207, w_096_215, w_096_235, w_096_248, w_096_283, w_096_296, w_096_303, w_096_330;
  wire w_097_008, w_097_025, w_097_027, w_097_036, w_097_064, w_097_067, w_097_070, w_097_092, w_097_097, w_097_111, w_097_114, w_097_125, w_097_133, w_097_139, w_097_146, w_097_148, w_097_163, w_097_164, w_097_165, w_097_167, w_097_182, w_097_188, w_097_193, w_097_205, w_097_215;
  wire w_098_004, w_098_005, w_098_006, w_098_008, w_098_009, w_098_010, w_098_011, w_098_013, w_098_014, w_098_015, w_098_016, w_098_017, w_098_018, w_098_020, w_098_022, w_098_023;
  wire w_099_006, w_099_013, w_099_015, w_099_020, w_099_022, w_099_026, w_099_037, w_099_038, w_099_043, w_099_052, w_099_054, w_099_056, w_099_059, w_099_075, w_099_088, w_099_110, w_099_111, w_099_120, w_099_123, w_099_150, w_099_159, w_099_164, w_099_180, w_099_181, w_099_196, w_099_223, w_099_226, w_099_244, w_099_267, w_099_271, w_099_277;
  wire w_100_003, w_100_035, w_100_041, w_100_046, w_100_062, w_100_127, w_100_149, w_100_157, w_100_163, w_100_179, w_100_180, w_100_193, w_100_194, w_100_215, w_100_219, w_100_230, w_100_231, w_100_258, w_100_273, w_100_298, w_100_301, w_100_312, w_100_402;
  wire w_101_001, w_101_002, w_101_010, w_101_015, w_101_019, w_101_023, w_101_024, w_101_030, w_101_034, w_101_039, w_101_043, w_101_048, w_101_052, w_101_054, w_101_065, w_101_074, w_101_078, w_101_099, w_101_101, w_101_105, w_101_106, w_101_126, w_101_128, w_101_145, w_101_158, w_101_163, w_101_175, w_101_186, w_101_201, w_101_225, w_101_249, w_101_254, w_101_270, w_101_301, w_101_305, w_101_329;
  wire w_102_003, w_102_013, w_102_028, w_102_030, w_102_031, w_102_036, w_102_039, w_102_044, w_102_047, w_102_059, w_102_071, w_102_076, w_102_077, w_102_078, w_102_079, w_102_080, w_102_083, w_102_087, w_102_094, w_102_097, w_102_111, w_102_127, w_102_129, w_102_131, w_102_147, w_102_149, w_102_155;
  wire w_103_000, w_103_001, w_103_002, w_103_003, w_103_004, w_103_005, w_103_006, w_103_007, w_103_008, w_103_009, w_103_011, w_103_012, w_103_013, w_103_015, w_103_016, w_103_017, w_103_018;
  wire w_104_002, w_104_007, w_104_014, w_104_022, w_104_026, w_104_031, w_104_034, w_104_045, w_104_061, w_104_112, w_104_129, w_104_192, w_104_223, w_104_260, w_104_263, w_104_301, w_104_303, w_104_327, w_104_365, w_104_373, w_104_374, w_104_379, w_104_385, w_104_430;
  wire w_105_001, w_105_012, w_105_026, w_105_033, w_105_035, w_105_041, w_105_047, w_105_051, w_105_057, w_105_077, w_105_078, w_105_116, w_105_121, w_105_123, w_105_129, w_105_151, w_105_165, w_105_167, w_105_177, w_105_192, w_105_231, w_105_246, w_105_248, w_105_293, w_105_297, w_105_317, w_105_382, w_105_426;
  wire w_106_003, w_106_007, w_106_010, w_106_022, w_106_079, w_106_109, w_106_146, w_106_164, w_106_168, w_106_176, w_106_184, w_106_202, w_106_211, w_106_232, w_106_262, w_106_269, w_106_271, w_106_286, w_106_295, w_106_337, w_106_342, w_106_354, w_106_359, w_106_380, w_106_395, w_106_408, w_106_422, w_106_482;
  wire w_107_003, w_107_010, w_107_013, w_107_021, w_107_022, w_107_023, w_107_032, w_107_040, w_107_041, w_107_043, w_107_045, w_107_046, w_107_047, w_107_056, w_107_057, w_107_058, w_107_061, w_107_067, w_107_068, w_107_069;
  wire w_108_000, w_108_008, w_108_010, w_108_011, w_108_017, w_108_019, w_108_023, w_108_024, w_108_025, w_108_028, w_108_029, w_108_030, w_108_032, w_108_036, w_108_038, w_108_040, w_108_043, w_108_045, w_108_046, w_108_050, w_108_056;
  wire w_109_000, w_109_001;
  wire w_110_005, w_110_007, w_110_008, w_110_020, w_110_027, w_110_034, w_110_035, w_110_041, w_110_049, w_110_051, w_110_060, w_110_094, w_110_095, w_110_132, w_110_142, w_110_149, w_110_156, w_110_161, w_110_172, w_110_193, w_110_194, w_110_210;
  wire w_111_001, w_111_005, w_111_007, w_111_014, w_111_015, w_111_017, w_111_020, w_111_024, w_111_028, w_111_030, w_111_036, w_111_037, w_111_047, w_111_048, w_111_055, w_111_061, w_111_066, w_111_069, w_111_081, w_111_087, w_111_088;
  wire w_112_017, w_112_020, w_112_028, w_112_033, w_112_035, w_112_050, w_112_053, w_112_071, w_112_073, w_112_074, w_112_078, w_112_081, w_112_098, w_112_103, w_112_105, w_112_108, w_112_131, w_112_142, w_112_150, w_112_156, w_112_184, w_112_212, w_112_232, w_112_304, w_112_363;
  wire w_113_002, w_113_007, w_113_010, w_113_014, w_113_020, w_113_030, w_113_035, w_113_039, w_113_041, w_113_042, w_113_045, w_113_048, w_113_052, w_113_056, w_113_059, w_113_062, w_113_066, w_113_072, w_113_075;
  wire w_114_001, w_114_015, w_114_022, w_114_027, w_114_038, w_114_040, w_114_048, w_114_050, w_114_057, w_114_058, w_114_077, w_114_080, w_114_092, w_114_098, w_114_102, w_114_115, w_114_146, w_114_153, w_114_159, w_114_181, w_114_187, w_114_188, w_114_192, w_114_195, w_114_208, w_114_237, w_114_266, w_114_267, w_114_268, w_114_269, w_114_270, w_114_271, w_114_272, w_114_273, w_114_274, w_114_275, w_114_276, w_114_278, w_114_280, w_114_281, w_114_282, w_114_283, w_114_284, w_114_285, w_114_286, w_114_287, w_114_289;
  wire w_115_031, w_115_032, w_115_037, w_115_095, w_115_131, w_115_164, w_115_171, w_115_174, w_115_185, w_115_195, w_115_203, w_115_212, w_115_242, w_115_247, w_115_308, w_115_314, w_115_320, w_115_330, w_115_346, w_115_379, w_115_423, w_115_424;
  wire w_116_022, w_116_023, w_116_026, w_116_028, w_116_029, w_116_037, w_116_038, w_116_054, w_116_059, w_116_094, w_116_100, w_116_108, w_116_116, w_116_137, w_116_191, w_116_202, w_116_208, w_116_214, w_116_218, w_116_243, w_116_275;
  wire w_117_016, w_117_060, w_117_138, w_117_157, w_117_161, w_117_176, w_117_201, w_117_221, w_117_238, w_117_261, w_117_266, w_117_279, w_117_289, w_117_294, w_117_322, w_117_324, w_117_325, w_117_341, w_117_344, w_117_353, w_117_357, w_117_362, w_117_375, w_117_386, w_117_403, w_117_406, w_117_410, w_117_411, w_117_414, w_117_434, w_117_449;
  wire w_118_020, w_118_024, w_118_026, w_118_046, w_118_054, w_118_060, w_118_080, w_118_084, w_118_104, w_118_108, w_118_141, w_118_172, w_118_175, w_118_187, w_118_194, w_118_196, w_118_217, w_118_242, w_118_277, w_118_293, w_118_297, w_118_310, w_118_329;
  wire w_119_001, w_119_006, w_119_040, w_119_101, w_119_107, w_119_114, w_119_122, w_119_136, w_119_141, w_119_157, w_119_168, w_119_184, w_119_187, w_119_222, w_119_250, w_119_279, w_119_282, w_119_287;
  wire w_120_004, w_120_009, w_120_016, w_120_021, w_120_040, w_120_043, w_120_045, w_120_061, w_120_063, w_120_064, w_120_065, w_120_070, w_120_086, w_120_088, w_120_089, w_120_092, w_120_109, w_120_110, w_120_115, w_120_117, w_120_136, w_120_140, w_120_168, w_120_193;
  wire w_121_001, w_121_034, w_121_035, w_121_054, w_121_070, w_121_090, w_121_096, w_121_107, w_121_126, w_121_128, w_121_159, w_121_164, w_121_242, w_121_247, w_121_269, w_121_284, w_121_300;
  wire w_122_002, w_122_004, w_122_014, w_122_021, w_122_026, w_122_028, w_122_034, w_122_045, w_122_057, w_122_079, w_122_084, w_122_086, w_122_089, w_122_092, w_122_096, w_122_107, w_122_110, w_122_113, w_122_114, w_122_125, w_122_128, w_122_141, w_122_152, w_122_157, w_122_161, w_122_163;
  wire w_123_007, w_123_012, w_123_023, w_123_026, w_123_030, w_123_055, w_123_062, w_123_067, w_123_068, w_123_075, w_123_077, w_123_078, w_123_082, w_123_087, w_123_120, w_123_124, w_123_149, w_123_167, w_123_188, w_123_210, w_123_255, w_123_265, w_123_296, w_123_326;
  wire w_124_001, w_124_002, w_124_020, w_124_030, w_124_031, w_124_078, w_124_088, w_124_099, w_124_106, w_124_116, w_124_147, w_124_162, w_124_174, w_124_211, w_124_234;
  wire w_125_010, w_125_030, w_125_081, w_125_117, w_125_132, w_125_152, w_125_165, w_125_166, w_125_186, w_125_222, w_125_234, w_125_239, w_125_246, w_125_249, w_125_255, w_125_359, w_125_396, w_125_411, w_125_463;
  wire w_126_001, w_126_005, w_126_009, w_126_012, w_126_016, w_126_020, w_126_024, w_126_036, w_126_040;
  wire w_127_016, w_127_021, w_127_033, w_127_075, w_127_133, w_127_140, w_127_172, w_127_189, w_127_237, w_127_246, w_127_256, w_127_260, w_127_272, w_127_328, w_127_368, w_127_371, w_127_404, w_127_492, w_127_493, w_127_494, w_127_495, w_127_496, w_127_497, w_127_498, w_127_499, w_127_500, w_127_501, w_127_502, w_127_503, w_127_505, w_127_507, w_127_508, w_127_509, w_127_510, w_127_511, w_127_512, w_127_513, w_127_514, w_127_515, w_127_516, w_127_517, w_127_519, w_127_521, w_127_522, w_127_523, w_127_524, w_127_525, w_127_526, w_127_527, w_127_528, w_127_529, w_127_530, w_127_531, w_127_532, w_127_534;
  wire w_128_013, w_128_015, w_128_025, w_128_031, w_128_032, w_128_034, w_128_038, w_128_042, w_128_043, w_128_045, w_128_048, w_128_051, w_128_054, w_128_057, w_128_058;
  wire w_129_000;
  wire w_130_009, w_130_012, w_130_021, w_130_027, w_130_034, w_130_037, w_130_068, w_130_072, w_130_086, w_130_087, w_130_106, w_130_107, w_130_111, w_130_137, w_130_142, w_130_146, w_130_171;
  wire w_131_001, w_131_009, w_131_012, w_131_024, w_131_040, w_131_041, w_131_058, w_131_063, w_131_081, w_131_127, w_131_141, w_131_142, w_131_169, w_131_191, w_131_196, w_131_198;
  wire w_132_037, w_132_054, w_132_067, w_132_100, w_132_104, w_132_113, w_132_114, w_132_133, w_132_169, w_132_176, w_132_182, w_132_185;
  wire w_133_026, w_133_068, w_133_076, w_133_101, w_133_174, w_133_227, w_133_232, w_133_282, w_133_357;
  wire w_134_002, w_134_003, w_134_004, w_134_020, w_134_022, w_134_026, w_134_033, w_134_034, w_134_042, w_134_043, w_134_046, w_134_047, w_134_053, w_134_054, w_134_062, w_134_063, w_134_064, w_134_068, w_134_069, w_134_073, w_134_075, w_134_085;
  wire w_135_027, w_135_049, w_135_097, w_135_113, w_135_115, w_135_123, w_135_131, w_135_153, w_135_186, w_135_203, w_135_222, w_135_250;
  wire w_136_001, w_136_002, w_136_007, w_136_013, w_136_014, w_136_017, w_136_018, w_136_019, w_136_021, w_136_022, w_136_029;
  wire w_137_008, w_137_010, w_137_014, w_137_021, w_137_031, w_137_035, w_137_041, w_137_045, w_137_050, w_137_054, w_137_057;
  wire w_138_006, w_138_013, w_138_122, w_138_128, w_138_174, w_138_215, w_138_217, w_138_223, w_138_241, w_138_242, w_138_243, w_138_244, w_138_245, w_138_246, w_138_247, w_138_248, w_138_252, w_138_253, w_138_254, w_138_255, w_138_256, w_138_257, w_138_259;
  wire w_139_016, w_139_025, w_139_030, w_139_043, w_139_112, w_139_150, w_139_154, w_139_164, w_139_176, w_139_182, w_139_187, w_139_188, w_139_229, w_139_230, w_139_231;
  wire w_140_005, w_140_026, w_140_043, w_140_044, w_140_049, w_140_071, w_140_080, w_140_084, w_140_106, w_140_110, w_140_157, w_140_196, w_140_266, w_140_300;
  wire w_141_005, w_141_022, w_141_061, w_141_122, w_141_153, w_141_154, w_141_163, w_141_169, w_141_172, w_141_193, w_141_207, w_141_261;
  wire w_142_000, w_142_070, w_142_078, w_142_083, w_142_086, w_142_098, w_142_103, w_142_106, w_142_111, w_142_116, w_142_122, w_142_131, w_142_146, w_142_150, w_142_173, w_142_176, w_142_204, w_142_250, w_142_279, w_142_303;
  wire w_143_002, w_143_018, w_143_025, w_143_033, w_143_054, w_143_061, w_143_070, w_143_087, w_143_088, w_143_092, w_143_099, w_143_103, w_143_107;
  wire w_144_004, w_144_010, w_144_016, w_144_045, w_144_058, w_144_062, w_144_064, w_144_095, w_144_105, w_144_107, w_144_124, w_144_136, w_144_151, w_144_172, w_144_186;
  wire w_145_006, w_145_009, w_145_063, w_145_072, w_145_073, w_145_143, w_145_196, w_145_215, w_145_219, w_145_250, w_145_333, w_145_393;
  wire w_146_011, w_146_017, w_146_033, w_146_037, w_146_041, w_146_050, w_146_061, w_146_064, w_146_087, w_146_161, w_146_168, w_146_200, w_146_220, w_146_228, w_146_245, w_146_307;
  wire w_147_012, w_147_019, w_147_033, w_147_063, w_147_066, w_147_074, w_147_084, w_147_106, w_147_107, w_147_119, w_147_127, w_147_129, w_147_136, w_147_138, w_147_151, w_147_175, w_147_191;
  wire w_148_012, w_148_022, w_148_028, w_148_038, w_148_069, w_148_073, w_148_087, w_148_121, w_148_129, w_148_242, w_148_251, w_148_324;
  wire w_149_000, w_149_001, w_149_003, w_149_004, w_149_005, w_149_007, w_149_008, w_149_011, w_149_018, w_149_019, w_149_022, w_149_023, w_149_024, w_149_026, w_149_027, w_149_028;
  wire w_150_024, w_150_063, w_150_082, w_150_089, w_150_106, w_150_122, w_150_146, w_150_156, w_150_176, w_150_225, w_150_320, w_150_334, w_150_392;
  wire w_151_000, w_151_007, w_151_008, w_151_010, w_151_021, w_151_023, w_151_029, w_151_033, w_151_034, w_151_036, w_151_038, w_151_041;
  wire w_152_022, w_152_029, w_152_032, w_152_050, w_152_053, w_152_056, w_152_059, w_152_062, w_152_072, w_152_083, w_152_120, w_152_132, w_152_134, w_152_147, w_152_191;
  wire w_153_001, w_153_007, w_153_008, w_153_025, w_153_093, w_153_108, w_153_125, w_153_186, w_153_209, w_153_218, w_153_255, w_153_297, w_153_331, w_153_409, w_153_424, w_153_461;
  wire w_154_009, w_154_013, w_154_024, w_154_047, w_154_050, w_154_051, w_154_058, w_154_062, w_154_075, w_154_078, w_154_103, w_154_106;
  wire w_155_023, w_155_072, w_155_080, w_155_101, w_155_102, w_155_110, w_155_165, w_155_189, w_155_231, w_155_237, w_155_261, w_155_272, w_155_322, w_155_329;
  wire w_156_066, w_156_090, w_156_115, w_156_144, w_156_153, w_156_168, w_156_217, w_156_225, w_156_302;
  wire w_157_019, w_157_165, w_157_229, w_157_242, w_157_393, w_157_434;
  wire w_158_000, w_158_001, w_158_003, w_158_006, w_158_007, w_158_011, w_158_013, w_158_016, w_158_025, w_158_027, w_158_036, w_158_038, w_158_039, w_158_040, w_158_041, w_158_042, w_158_043, w_158_044, w_158_045, w_158_046, w_158_047, w_158_048;
  wire w_159_005, w_159_007, w_159_055, w_159_072, w_159_073, w_159_080, w_159_092, w_159_107, w_159_128, w_159_158, w_159_199, w_159_210;
  wire w_160_013, w_160_014, w_160_025, w_160_060, w_160_071, w_160_072, w_160_075, w_160_102, w_160_114, w_160_132, w_160_138;
  wire w_161_013, w_161_031, w_161_039, w_161_067, w_161_083, w_161_141, w_161_153, w_161_160, w_161_171, w_161_207, w_161_219, w_161_261;
  wire w_162_000, w_162_001, w_162_005, w_162_007, w_162_008, w_162_009, w_162_010, w_162_011, w_162_012, w_162_013, w_162_014, w_162_015, w_162_017;
  wire w_163_000, w_163_003, w_163_007, w_163_016, w_163_035, w_163_054, w_163_070, w_163_133, w_163_147, w_163_156, w_163_171, w_163_187, w_163_210, w_163_250, w_163_330, w_163_371, w_163_383;
  wire w_164_001, w_164_012, w_164_020, w_164_027, w_164_058, w_164_090, w_164_098, w_164_106, w_164_119, w_164_132, w_164_136, w_164_163, w_164_188, w_164_189, w_164_190, w_164_191, w_164_192, w_164_193, w_164_194, w_164_195;
  wire w_165_004, w_165_028, w_165_057, w_165_092, w_165_104, w_165_111, w_165_112, w_165_174, w_165_282, w_165_293, w_165_339;
  wire w_166_021, w_166_042, w_166_075, w_166_112, w_166_181, w_166_250, w_166_255;
  wire w_167_011, w_167_035, w_167_037, w_167_053, w_167_109, w_167_136, w_167_138, w_167_152, w_167_157, w_167_168, w_167_231, w_167_302;
  wire w_168_002, w_168_011, w_168_015, w_168_046, w_168_047, w_168_053, w_168_054, w_168_082, w_168_103, w_168_115, w_168_138, w_168_143, w_168_145, w_168_151, w_168_157;
  wire w_169_072, w_169_215, w_169_216, w_169_217, w_169_222;
  wire w_170_029, w_170_038, w_170_061, w_170_083, w_170_089, w_170_098, w_170_112, w_170_137, w_170_145, w_170_175, w_170_190, w_170_198, w_170_216, w_170_219, w_170_221, w_170_248;
  wire w_171_029, w_171_084, w_171_110, w_171_121, w_171_152, w_171_173, w_171_227, w_171_268, w_171_276;
  wire w_172_009, w_172_012, w_172_018, w_172_041, w_172_052, w_172_094, w_172_102, w_172_111, w_172_152, w_172_168, w_172_207, w_172_224;
  wire w_173_003, w_173_004, w_173_062, w_173_086, w_173_101, w_173_121, w_173_134, w_173_145, w_173_204, w_173_206, w_173_209, w_173_221, w_173_267, w_173_271, w_173_283, w_173_284, w_173_285, w_173_286, w_173_287, w_173_288, w_173_289, w_173_290, w_173_291, w_173_292;
  wire w_174_063, w_174_090, w_174_144, w_174_147, w_174_209, w_174_253, w_174_278, w_174_323, w_174_378, w_174_399, w_174_416, w_174_492;
  wire w_175_045, w_175_077, w_175_099, w_175_137, w_175_171, w_175_173, w_175_203, w_175_214, w_175_262, w_175_274, w_175_373;
  wire w_176_036, w_176_067, w_176_095, w_176_111, w_176_144, w_176_196, w_176_240, w_176_242, w_176_372, w_176_380, w_176_383, w_176_396, w_176_397;
  wire w_177_001, w_177_043, w_177_089, w_177_152, w_177_212, w_177_215, w_177_222;
  wire w_178_029, w_178_049, w_178_080, w_178_104, w_178_121, w_178_172, w_178_304, w_178_334;
  wire w_179_002, w_179_084, w_179_138;
  wire w_180_007, w_180_013, w_180_070, w_180_120, w_180_133, w_180_178, w_180_204, w_180_208, w_180_210, w_180_279;
  wire w_181_041, w_181_047, w_181_056, w_181_066, w_181_073, w_181_082, w_181_087, w_181_089, w_181_107, w_181_119;
  wire w_182_000, w_182_004, w_182_010, w_182_016, w_182_021, w_182_024, w_182_026, w_182_033, w_182_035, w_182_039, w_182_046, w_182_059, w_182_077, w_182_080, w_182_087, w_182_094, w_182_100;
  wire w_183_019, w_183_036, w_183_038, w_183_077;
  wire w_184_015, w_184_021, w_184_056, w_184_069, w_184_095, w_184_139, w_184_158, w_184_178, w_184_185, w_184_246, w_184_289, w_184_368, w_184_393, w_184_412, w_184_418, w_184_450;
  wire w_185_031, w_185_076, w_185_109, w_185_122, w_185_123, w_185_126, w_185_270;
  wire w_186_008, w_186_024, w_186_038, w_186_052, w_186_053, w_186_056, w_186_061, w_186_062, w_186_063, w_186_064, w_186_065, w_186_066, w_186_067, w_186_068, w_186_072, w_186_073, w_186_074, w_186_075, w_186_076, w_186_077, w_186_078, w_186_079, w_186_080, w_186_081, w_186_082, w_186_083, w_186_085;
  wire w_187_032, w_187_053, w_187_131, w_187_155, w_187_159;
  wire w_188_011, w_188_034, w_188_047, w_188_048, w_188_081, w_188_089, w_188_101, w_188_105, w_188_109;
  wire w_189_029, w_189_058, w_189_062, w_189_067, w_189_135, w_189_145, w_189_213, w_189_303;
  wire w_190_014, w_190_015, w_190_025, w_190_027, w_190_042, w_190_066, w_190_077, w_190_081, w_190_102;
  wire w_191_004, w_191_024, w_191_075, w_191_082, w_191_092, w_191_150, w_191_156, w_191_174, w_191_181;
  wire w_192_024, w_192_062, w_192_086, w_192_129, w_192_206, w_192_221, w_192_230, w_192_247, w_192_260, w_192_261, w_192_262, w_192_263, w_192_264, w_192_265, w_192_266, w_192_267, w_192_268;
  wire w_193_012, w_193_023, w_193_039, w_193_048, w_193_082;
  wire w_194_013, w_194_058, w_194_252, w_194_259, w_194_273;
  wire w_195_016, w_195_041, w_195_053, w_195_058, w_195_061, w_195_076, w_195_080, w_195_081, w_195_082;
  wire w_196_023, w_196_069, w_196_070, w_196_096, w_196_141, w_196_211, w_196_214, w_196_245, w_196_247;
  wire w_197_024, w_197_033, w_197_081, w_197_083, w_197_098, w_197_102, w_197_103, w_197_142, w_197_174, w_197_206;
  wire w_198_020, w_198_030, w_198_071, w_198_093, w_198_111, w_198_179, w_198_225, w_198_323, w_198_338, w_198_350;
  wire w_199_006, w_199_007, w_199_014, w_199_018, w_199_019, w_199_021, w_199_026;
  wire w_200_011, w_200_025, w_200_028, w_200_085, w_200_130, w_200_186, w_200_204, w_200_235, w_200_253, w_200_254;
  wire w_201_007, w_201_017, w_201_024, w_201_039, w_201_090, w_201_127, w_201_196, w_201_204, w_201_344;
  wire w_202_032, w_202_056, w_202_150, w_202_207, w_202_230, w_202_303, w_202_311, w_202_411, w_202_416;
  wire w_203_038, w_203_055, w_203_066, w_203_071, w_203_093, w_203_235, w_203_367, w_203_368, w_203_369, w_203_370, w_203_371, w_203_372, w_203_373, w_203_377, w_203_378, w_203_379, w_203_380, w_203_381, w_203_382, w_203_383, w_203_384, w_203_385, w_203_386, w_203_387, w_203_388, w_203_390;
  wire w_204_014, w_204_034, w_204_058, w_204_066, w_204_083, w_204_117, w_204_135, w_204_223, w_204_239, w_204_260, w_204_274;
  wire w_205_004, w_205_007, w_205_023, w_205_047, w_205_051, w_205_066;
  wire w_206_030, w_206_035, w_206_063, w_206_098, w_206_162, w_206_222, w_206_238, w_206_331;
  wire w_207_027, w_207_041, w_207_130, w_207_204, w_207_277, w_207_303;
  wire w_208_001, w_208_004, w_208_022, w_208_024, w_208_032, w_208_037, w_208_052, w_208_076, w_208_086, w_208_126;
  wire w_209_033, w_209_063, w_209_080, w_209_129, w_209_148, w_209_406;
  wire w_210_032, w_210_060, w_210_136, w_210_140, w_210_164, w_210_167, w_210_176, w_210_212, w_210_213, w_210_216, w_210_226, w_210_228;
  wire w_211_055, w_211_058, w_211_075, w_211_077, w_211_095, w_211_118, w_211_135, w_211_136, w_211_257;
  wire w_212_031, w_212_037, w_212_052, w_212_054, w_212_063, w_212_123, w_212_172, w_212_192;
  wire w_213_007, w_213_014, w_213_044, w_213_071, w_213_177;
  wire w_214_020, w_214_023, w_214_026, w_214_029, w_214_039, w_214_047, w_214_053, w_214_054, w_214_056;
  wire w_215_008, w_215_035, w_215_054, w_215_063, w_215_075, w_215_085, w_215_102, w_215_170, w_215_221, w_215_228, w_215_234;
  wire w_216_003, w_216_017, w_216_041, w_216_050, w_216_067, w_216_072, w_216_076, w_216_123;
  wire w_217_088, w_217_326, w_217_420, w_217_423, w_217_434;
  wire w_218_031, w_218_048, w_218_068, w_218_081, w_218_163, w_218_287, w_218_396;
  wire w_219_011, w_219_041, w_219_086, w_219_220, w_219_246, w_219_254, w_219_260, w_219_263, w_219_290, w_219_300, w_219_314, w_219_361;
  wire w_220_054, w_220_254, w_220_258, w_220_261, w_220_315, w_220_358, w_220_440, w_220_449, w_220_480;
  wire w_221_012, w_221_046, w_221_050, w_221_064, w_221_079, w_221_099, w_221_102, w_221_107, w_221_113;
  wire w_222_028, w_222_030, w_222_067, w_222_086, w_222_100, w_222_218, w_222_264;
  wire w_223_066, w_223_074, w_223_095, w_223_099, w_223_168, w_223_194;
  wire w_224_000, w_224_001, w_224_012, w_224_016, w_224_017, w_224_038, w_224_045, w_224_053;
  wire w_225_005, w_225_059, w_225_069, w_225_167, w_225_184, w_225_224, w_225_248;
  wire w_226_101, w_226_153, w_226_188, w_226_202, w_226_310, w_226_336, w_226_396, w_226_397, w_226_398, w_226_399, w_226_400, w_226_401, w_226_402, w_226_403;
  wire w_227_019, w_227_038, w_227_059, w_227_061, w_227_076, w_227_112, w_227_150, w_227_218, w_227_243, w_227_285, w_227_330;
  wire w_228_041, w_228_066, w_228_087, w_228_098, w_228_284;
  wire w_229_058, w_229_092, w_229_140, w_229_181, w_229_269;
  wire w_230_013, w_230_017, w_230_025, w_230_036, w_230_043, w_230_053, w_230_054;
  wire w_231_000, w_231_005, w_231_041, w_231_046, w_231_049, w_231_064, w_231_066;
  wire w_232_075;
  wire w_233_031, w_233_065, w_233_083, w_233_104, w_233_203, w_233_305;
  wire w_234_001, w_234_093, w_234_099, w_234_115, w_234_117, w_234_122;
  wire w_235_118, w_235_211;
  wire w_236_005, w_236_011, w_236_018, w_236_024, w_236_027, w_236_043, w_236_046, w_236_068;
  wire w_237_008, w_237_011, w_237_025, w_237_037;
  wire w_238_043, w_238_092, w_238_094, w_238_126, w_238_130, w_238_170, w_238_190, w_238_262, w_238_272, w_238_309, w_238_319;
  wire w_239_017, w_239_061, w_239_068, w_239_092, w_239_096, w_239_152, w_239_236, w_239_311;
  wire w_240_026, w_240_041, w_240_046, w_240_072, w_240_122, w_240_180, w_240_182, w_240_196, w_240_206, w_240_213;
  wire w_241_014, w_241_017, w_241_021, w_241_047, w_241_053, w_241_074;
  wire w_242_038, w_242_105, w_242_163, w_242_346;
  wire w_243_190;
  wire w_244_022, w_244_075, w_244_089, w_244_109, w_244_135, w_244_160;
  wire w_245_019, w_245_057, w_245_106, w_245_118, w_245_121, w_245_135, w_245_193;
  wire w_246_019, w_246_065, w_246_078, w_246_093, w_246_258, w_246_273, w_246_363;
  wire w_247_040, w_247_054, w_247_065, w_247_223, w_247_230, w_247_254;
  wire w_248_029, w_248_115, w_248_133, w_248_243, w_248_360;
  wire w_249_029, w_249_031, w_249_033, w_249_052, w_249_068, w_249_082, w_249_083, w_249_089, w_249_102;
  wire w_250_002, w_250_029, w_250_035, w_250_044, w_250_047, w_250_049, w_250_057;
  wire w_251_017, w_251_038, w_251_056, w_251_085, w_251_098, w_251_112, w_251_113, w_251_124;
  wire w_252_002, w_252_041, w_252_092, w_252_147, w_252_234, w_252_279, w_252_327, w_252_383;
  wire w_253_010, w_253_023, w_253_048, w_253_097, w_253_123, w_253_140;
  wire w_254_014, w_254_037, w_254_050, w_254_101;
  wire w_255_037, w_255_057, w_255_068, w_255_186, w_255_197;
  wire w_256_005, w_256_011, w_256_072, w_256_125, w_256_134;
  wire w_257_014, w_257_040, w_257_048, w_257_050, w_257_052, w_257_073, w_257_102, w_257_168, w_257_213, w_257_214;
  wire w_258_022, w_258_045, w_258_046, w_258_190, w_258_261;
  wire w_259_042, w_259_044, w_259_079, w_259_102, w_259_104, w_259_131, w_259_153;
  wire w_260_000, w_260_054, w_260_057, w_260_063, w_260_074, w_260_076, w_260_163, w_260_181;
  wire w_261_041, w_261_083, w_261_115;
  wire w_262_050, w_262_063, w_262_064, w_262_065, w_262_066, w_262_067, w_262_068, w_262_069, w_262_070, w_262_071, w_262_072, w_262_073, w_262_074;
  wire w_263_020, w_263_026, w_263_040, w_263_053, w_263_114, w_263_194;
  wire w_264_012, w_264_064, w_264_085, w_264_125, w_264_191, w_264_275, w_264_355;
  wire w_265_000, w_265_003, w_265_006, w_265_017;
  wire w_266_076, w_266_111, w_266_314, w_266_408;
  wire w_267_128, w_267_222, w_267_355, w_267_389;
  wire w_268_018, w_268_025, w_268_040, w_268_139, w_268_150;
  wire w_269_029, w_269_038, w_269_043, w_269_055, w_269_059;
  wire w_270_021, w_270_054, w_270_111, w_270_190, w_270_255;
  wire w_271_026, w_271_048, w_271_118, w_271_151, w_271_172, w_271_254, w_271_280, w_271_338;
  wire w_272_003, w_272_009, w_272_010, w_272_019, w_272_020, w_272_022, w_272_024, w_272_029, w_272_031;
  wire w_273_023, w_273_044, w_273_071, w_273_142, w_273_143;
  wire w_274_017, w_274_034, w_274_149, w_274_192;
  wire w_275_053, w_275_054, w_275_088, w_275_097, w_275_117, w_275_123;
  wire w_276_117;
  wire w_277_003, w_277_005, w_277_013, w_277_015, w_277_046;
  wire w_278_079, w_278_118;
  wire w_279_071, w_279_309, w_279_345, w_279_415;
  wire w_280_008, w_280_025, w_280_060, w_280_063;
  wire w_281_002, w_281_009, w_281_010, w_281_015, w_281_016;
  wire w_282_037, w_282_046, w_282_065, w_282_096, w_282_122;
  wire w_283_026, w_283_139, w_283_169, w_283_188, w_283_224;
  wire w_284_013, w_284_122, w_284_265;
  wire w_285_000, w_285_018, w_285_021, w_285_022, w_285_025, w_285_026, w_285_027, w_285_028, w_285_029, w_285_030, w_285_031, w_285_032, w_285_033, w_285_034, w_285_035;
  wire w_286_002, w_286_039, w_286_054, w_286_088, w_286_234, w_286_434;
  wire w_287_000, w_287_135, w_287_179, w_287_254, w_287_256, w_287_308, w_287_423, w_287_477;
  wire w_288_027, w_288_190;
  wire w_289_079, w_289_089, w_289_097, w_289_099, w_289_118, w_289_120, w_289_124;
  wire w_290_019, w_290_069;
  wire w_291_015, w_291_122, w_291_131;
  wire w_292_087, w_292_099, w_292_106;
  wire w_293_011, w_293_037, w_293_099, w_293_134;
  wire w_294_001, w_294_037, w_294_111, w_294_185;
  wire w_295_050, w_295_090, w_295_171, w_295_208, w_295_315;
  wire w_296_135, w_296_144, w_296_401, w_296_411;
  wire w_297_016, w_297_021, w_297_027, w_297_038, w_297_287, w_297_365;
  wire w_298_024, w_298_031, w_298_112, w_298_179, w_298_191;
  wire w_299_032;
  wire w_300_121, w_300_202, w_300_233, w_300_250;
  wire w_301_027, w_301_161;
  wire w_302_029, w_302_079, w_302_097, w_302_103;
  wire w_303_011, w_303_084, w_303_127, w_303_144, w_303_162, w_303_178, w_303_197, w_303_198, w_303_199, w_303_200, w_303_204, w_303_205, w_303_206, w_303_207, w_303_208, w_303_209, w_303_210, w_303_211, w_303_212, w_303_213, w_303_215;
  wire w_304_065, w_304_136, w_304_188;
  wire w_305_007, w_305_054, w_305_057, w_305_085;
  wire w_306_004, w_306_007, w_306_088, w_306_287;
  wire w_307_002, w_307_062, w_307_075, w_307_123, w_307_129, w_307_183;
  wire w_308_024, w_308_027, w_308_050;
  wire w_309_026, w_309_065, w_309_073, w_309_095, w_309_115, w_309_145;
  wire w_310_070, w_310_071, w_310_072, w_310_184, w_310_226;
  wire w_311_067, w_311_134, w_311_149, w_311_174;
  wire w_312_068, w_312_123, w_312_137, w_312_171, w_312_174, w_312_199, w_312_222;
  wire w_313_074, w_313_089, w_313_092, w_313_111, w_313_119, w_313_151;
  wire w_314_093, w_314_142, w_314_214, w_314_369, w_314_382;
  wire w_315_122, w_315_242, w_315_288, w_315_325;
  wire w_316_014, w_316_021, w_316_044, w_316_046, w_316_057, w_316_224;
  wire w_317_116, w_317_248, w_317_304, w_317_341, w_317_342, w_317_343, w_317_344, w_317_345, w_317_346, w_317_347, w_317_348, w_317_349, w_317_350, w_317_351;
  wire w_318_049, w_318_084, w_318_159, w_318_290, w_318_309, w_318_342, w_318_382, w_318_383, w_318_384, w_318_385, w_318_386, w_318_387, w_318_388, w_318_389, w_318_390, w_318_394, w_318_395, w_318_396, w_318_397, w_318_398, w_318_399, w_318_401;
  wire w_319_007, w_319_030, w_319_064, w_319_081, w_319_099;
  wire w_320_108, w_320_219, w_320_260;
  wire w_321_001, w_321_056, w_321_096, w_321_108;
  wire w_322_007, w_322_030;
  wire w_323_000, w_323_003, w_323_033, w_323_046, w_323_057;
  wire w_324_047;
  wire w_325_126, w_325_190, w_325_206, w_325_464;
  wire w_326_028, w_326_035, w_326_040, w_326_053, w_326_069;
  wire w_327_041, w_327_163, w_327_172, w_327_176;
  wire w_328_038, w_328_058, w_328_215, w_328_241, w_328_297, w_328_459;
  wire w_329_074, w_329_237, w_329_287, w_329_321, w_329_342, w_329_431;
  wire w_330_029, w_330_134, w_330_154, w_330_364;
  wire w_331_017, w_331_022, w_331_032, w_331_042;
  wire w_332_014, w_332_197, w_332_226, w_332_255;
  wire w_333_072, w_333_074, w_333_091, w_333_179;
  wire w_334_478;
  wire w_335_029, w_335_044, w_335_066, w_335_091, w_335_121, w_335_209;
  wire w_336_060, w_336_091, w_336_289, w_336_307;
  wire w_337_030, w_337_118, w_337_195, w_337_215;
  wire w_338_026, w_338_063, w_338_069, w_338_278, w_338_330, w_338_357, w_338_358, w_338_359, w_338_360, w_338_361, w_338_362;
  wire w_339_007, w_339_051, w_339_053, w_339_177;
  wire w_340_000, w_340_011, w_340_014, w_340_040, w_340_054, w_340_055, w_340_057, w_340_109;
  wire w_341_000;
  wire w_342_008, w_342_045, w_342_047, w_342_126, w_342_127;
  wire w_343_007, w_343_037, w_343_039, w_343_135, w_343_174, w_343_228, w_343_266;
  wire w_344_173, w_344_199, w_344_457;
  wire w_345_011, w_345_135, w_345_273, w_345_274;
  wire w_346_050, w_346_109, w_346_129, w_346_130, w_346_227;
  wire w_347_016, w_347_336;
  wire w_348_014, w_348_030, w_348_081;
  wire w_349_191, w_349_245, w_349_281;
  wire w_350_004, w_350_028, w_350_047, w_350_238;
  wire w_351_071, w_351_146, w_351_203, w_351_242;
  wire w_353_014, w_353_076, w_353_085, w_353_130;
  wire w_354_003, w_354_039, w_354_041, w_354_079;
  wire w_355_015, w_355_017, w_355_028;
  wire w_356_143, w_356_161;
  wire w_357_008, w_357_130, w_357_180;
  wire w_358_387, w_358_405;
  wire w_359_035, w_359_038;
  wire w_360_045, w_360_064, w_360_083, w_360_088, w_360_148, w_360_183;
  wire w_361_066, w_361_099;
  wire w_362_046, w_362_069;
  wire w_363_010, w_363_018, w_363_068, w_363_072, w_363_094, w_363_100;
  wire w_364_037, w_364_083, w_364_094, w_364_121, w_364_172, w_364_241, w_364_268;
  wire w_365_028, w_365_042, w_365_077, w_365_141;
  wire w_366_026, w_366_124, w_366_148, w_366_183, w_366_193, w_366_206;
  wire w_367_049, w_367_165, w_367_393;
  wire w_368_097, w_368_099;
  wire w_369_179, w_369_376;
  wire w_370_025, w_370_064, w_370_123, w_370_137;
  wire w_371_122, w_371_325;
  wire w_372_024, w_372_062, w_372_070, w_372_147, w_372_148, w_372_149, w_372_150, w_372_151, w_372_152, w_372_153, w_372_154;
  wire w_373_007, w_373_024, w_373_071, w_373_092, w_373_093, w_373_102, w_373_103, w_373_104, w_373_105, w_373_106, w_373_107;
  wire w_374_002, w_374_034, w_374_035, w_374_110;
  wire w_375_169, w_375_263, w_375_264, w_375_265, w_375_266, w_375_267, w_375_268, w_375_269, w_375_270, w_375_271, w_375_272, w_375_276, w_375_277, w_375_278, w_375_279, w_375_280, w_375_281, w_375_282, w_375_283, w_375_284, w_375_285, w_375_286, w_375_288;
  wire w_376_092, w_376_151;
  wire w_377_008, w_377_053, w_377_379;
  wire w_378_049, w_378_126, w_378_141, w_378_179;
  wire w_379_118;
  wire w_380_152, w_380_293, w_380_334;
  wire w_381_074, w_381_248, w_381_443;
  wire w_382_002, w_382_034, w_382_056;
  wire w_383_159;
  wire w_384_042, w_384_057, w_384_072;
  wire w_385_013, w_385_014, w_385_064;
  wire w_386_035, w_386_178, w_386_290;
  wire w_387_024, w_387_051, w_387_113;
  wire w_388_115;
  wire w_389_033, w_389_067;
  wire w_390_001, w_390_052;
  wire w_392_137, w_392_288;
  wire w_393_155;
  wire w_394_016, w_394_020, w_394_024, w_394_050;
  wire w_395_002, w_395_203;
  wire w_396_016;
  wire w_398_176;
  wire w_399_000, w_399_010, w_399_015, w_399_028, w_399_043, w_399_049, w_399_054;
  wire w_400_010, w_400_042, w_400_047, w_400_075, w_400_084, w_400_091;
  wire w_401_091, w_401_410;
  wire w_402_009, w_402_035, w_402_045;
  wire w_403_036;
  wire w_404_279, w_404_377;
  wire w_405_041, w_405_167, w_405_178;
  wire w_407_015, w_407_108, w_407_159;
  wire w_408_002, w_408_030, w_408_171, w_408_216, w_408_271;
  wire w_409_254, w_409_279, w_409_310;
  wire w_410_005, w_410_075;
  wire w_411_149;
  wire w_412_009, w_412_010, w_412_014, w_412_037;
  wire w_413_022, w_413_029, w_413_052, w_413_064;
  wire w_414_028;
  wire w_415_029, w_415_041, w_415_054;
  wire w_416_296, w_416_319, w_416_450;
  wire w_417_006, w_417_038, w_417_103, w_417_133;
  wire w_418_069, w_418_107, w_418_144;
  wire w_419_064;
  wire w_420_044, w_420_081;
  wire w_421_002, w_421_026, w_421_038, w_421_047, w_421_048, w_421_063;
  wire w_423_034, w_423_087, w_423_090, w_423_096;
  wire w_424_100;
  wire w_425_154, w_425_195;
  wire w_426_047, w_426_084;
  wire w_427_195;
  wire w_428_147, w_428_176, w_428_202;
  wire w_429_028, w_429_123, w_429_342;
  wire w_430_100, w_430_237, w_430_283;
  wire w_431_065, w_431_155, w_431_274, w_431_275, w_431_276, w_431_277, w_431_281, w_431_282, w_431_283, w_431_284, w_431_285, w_431_286, w_431_287, w_431_288, w_431_290;
  wire w_432_071, w_432_131, w_432_234;
  wire w_433_039, w_433_297;
  wire w_434_098, w_434_174;
  wire w_436_036, w_436_131;
  wire w_437_142, w_437_314, w_437_372, w_437_387, w_437_409;
  wire w_438_037;
  wire w_439_040, w_439_186, w_439_302, w_439_333;
  wire w_440_021, w_440_090;
  wire w_441_005, w_441_048, w_441_160, w_441_164;
  wire w_442_039;
  wire w_443_013, w_443_224;
  wire w_444_092, w_444_099, w_444_139;
  wire w_445_002, w_445_239, w_445_354, w_445_400, w_445_401, w_445_402, w_445_403, w_445_404, w_445_408, w_445_409, w_445_410, w_445_411, w_445_412, w_445_413, w_445_414, w_445_416;
  wire w_446_008;
  wire w_447_052;
  wire w_448_017;
  wire w_450_061, w_450_294;
  wire w_452_024, w_452_134;
  wire w_453_014, w_453_051, w_453_349;
  wire w_454_080, w_454_088, w_454_409;
  wire w_455_005, w_455_008, w_455_023;
  wire w_456_263, w_456_272, w_456_397;
  wire w_458_002;
  wire w_459_250;
  wire w_460_219;
  wire w_461_097;
  wire w_462_065;
  wire w_463_068, w_463_096;
  wire w_464_100, w_464_175;
  wire w_465_019;
  wire w_467_079, w_467_208, w_467_415;
  wire w_468_311, w_468_341, w_468_377;
  wire w_469_026, w_469_317, w_469_331;
  wire w_471_034, w_471_092;
  wire w_472_120;
  wire w_473_338;
  wire w_474_062, w_474_179, w_474_313;
  wire w_475_091, w_475_104, w_475_130;
  wire w_476_067, w_476_252, w_476_253, w_476_254, w_476_255, w_476_256, w_476_257, w_476_258, w_476_259, w_476_260;
  wire w_477_036, w_477_047;
  wire w_478_218, w_478_276;
  wire w_479_094;
  wire w_480_000, w_480_002, w_480_004, w_480_008, w_480_010;
  wire w_481_017, w_481_077;
  wire w_482_000, w_482_001, w_482_008;
  wire w_483_015, w_483_041;
  wire w_484_029, w_484_092, w_484_093, w_484_094, w_484_095, w_484_096, w_484_100, w_484_101, w_484_102, w_484_103, w_484_105;
  wire w_485_027, w_485_084;
  wire w_486_007;
  wire w_487_030, w_487_053, w_487_054, w_487_064, w_487_077, w_487_078, w_487_079, w_487_083, w_487_084, w_487_085, w_487_086, w_487_087, w_487_088, w_487_089, w_487_090, w_487_091, w_487_092, w_487_093, w_487_094, w_487_096;
  wire w_488_206;
  wire w_489_323, w_489_324, w_489_325, w_489_326, w_489_327, w_489_328, w_489_329, w_489_330, w_489_331, w_489_332, w_489_336, w_489_337, w_489_338, w_489_339, w_489_340, w_489_341, w_489_342, w_489_344;
  wire w_490_000, w_490_172;
  wire w_492_089;
  wire w_498_010;
  wire w_500_000, w_500_001, w_500_002, w_500_003, w_500_004, w_500_005, w_500_006, w_500_007, w_500_008, w_500_009, w_500_010, w_500_011, w_500_012, w_500_013, w_500_014, w_500_015, w_500_016, w_500_017, w_500_018, w_500_019, w_500_020, w_500_021, w_500_022, w_500_023, w_500_024, w_500_025, w_500_026, w_500_027, w_500_028, w_500_029, w_500_030, w_500_031, w_500_032, w_500_033, w_500_034, w_500_035, w_500_036, w_500_037, w_500_038, w_500_039, w_500_040, w_500_041, w_500_042, w_500_043, w_500_044, w_500_045, w_500_046, w_500_047, w_500_048, w_500_049, w_500_050, w_500_051, w_500_052, w_500_053, w_500_054, w_500_055, w_500_056, w_500_057, w_500_058, w_500_059, w_500_060, w_500_061, w_500_062, w_500_063, w_500_064, w_500_065, w_500_066, w_500_067, w_500_068, w_500_069, w_500_070, w_500_071, w_500_072, w_500_073, w_500_074, w_500_075, w_500_076, w_500_077, w_500_078, w_500_079, w_500_080, w_500_081, w_500_082, w_500_083, w_500_084, w_500_085, w_500_086, w_500_087, w_500_088, w_500_089, w_500_090, w_500_091, w_500_092, w_500_093, w_500_094, w_500_095, w_500_096, w_500_097, w_500_098, w_500_099, w_500_100, w_500_101, w_500_102, w_500_103, w_500_104, w_500_105, w_500_106, w_500_107, w_500_108, w_500_109, w_500_110, w_500_111, w_500_112, w_500_113, w_500_114, w_500_115, w_500_116, w_500_117, w_500_118, w_500_119, w_500_120, w_500_121, w_500_122, w_500_123, w_500_124, w_500_125, w_500_126, w_500_127, w_500_128, w_500_129, w_500_130, w_500_131, w_500_132, w_500_133, w_500_134, w_500_135, w_500_136, w_500_137, w_500_138, w_500_139, w_500_140, w_500_141, w_500_142, w_500_143, w_500_144, w_500_145, w_500_146, w_500_147, w_500_148, w_500_149, w_500_150, w_500_151, w_500_152, w_500_153, w_500_154, w_500_155, w_500_156, w_500_157, w_500_158, w_500_159, w_500_160, w_500_161, w_500_162, w_500_163, w_500_164, w_500_165, w_500_166, w_500_167, w_500_168, w_500_169, w_500_170, w_500_171, w_500_172, w_500_173, w_500_174, w_500_175, w_500_176, w_500_177, w_500_178, w_500_179, w_500_180, w_500_181, w_500_182, w_500_183, w_500_184, w_500_185, w_500_186, w_500_187, w_500_188, w_500_189, w_500_190, w_500_191, w_500_192, w_500_193, w_500_194, w_500_195, w_500_196, w_500_197, w_500_198, w_500_199, w_500_200, w_500_201, w_500_202, w_500_203, w_500_204, w_500_205, w_500_206, w_500_207, w_500_208, w_500_209, w_500_210, w_500_211, w_500_212, w_500_213, w_500_214, w_500_215, w_500_216, w_500_217, w_500_218, w_500_219, w_500_220, w_500_221, w_500_222, w_500_223, w_500_224, w_500_225, w_500_226, w_500_227, w_500_228, w_500_229, w_500_230, w_500_231, w_500_232, w_500_233, w_500_234, w_500_235, w_500_236, w_500_237, w_500_238, w_500_239, w_500_240, w_500_241, w_500_242, w_500_243, w_500_244, w_500_245, w_500_246, w_500_247, w_500_248, w_500_249, w_500_250, w_500_251, w_500_252, w_500_253, w_500_254, w_500_255, w_500_256, w_500_257, w_500_258, w_500_259, w_500_260, w_500_261, w_500_262, w_500_263, w_500_264, w_500_265, w_500_266, w_500_267, w_500_268, w_500_269, w_500_270, w_500_271, w_500_272, w_500_273, w_500_274, w_500_275, w_500_276, w_500_277, w_500_278, w_500_279, w_500_280, w_500_281, w_500_282, w_500_283, w_500_284, w_500_285, w_500_286, w_500_287, w_500_288, w_500_289, w_500_290, w_500_291, w_500_292, w_500_293, w_500_294, w_500_295, w_500_296, w_500_297, w_500_298, w_500_299, w_500_300, w_500_301, w_500_302, w_500_303, w_500_304, w_500_305, w_500_306, w_500_307, w_500_308, w_500_309, w_500_310, w_500_311, w_500_312, w_500_313, w_500_314, w_500_315, w_500_316, w_500_317, w_500_318, w_500_319, w_500_320, w_500_321, w_500_322, w_500_323, w_500_324, w_500_325, w_500_326, w_500_327, w_500_328, w_500_329, w_500_330, w_500_331, w_500_332, w_500_333, w_500_334, w_500_335, w_500_336, w_500_337, w_500_338, w_500_339, w_500_340, w_500_341, w_500_342, w_500_343, w_500_344, w_500_345, w_500_346, w_500_347, w_500_348, w_500_349, w_500_350, w_500_351, w_500_352, w_500_353, w_500_354, w_500_355, w_500_356, w_500_357, w_500_358, w_500_359, w_500_360, w_500_361, w_500_362, w_500_363, w_500_364, w_500_365, w_500_366, w_500_367, w_500_368, w_500_369, w_500_370, w_500_371, w_500_372, w_500_373, w_500_374, w_500_375, w_500_376, w_500_377, w_500_378, w_500_379, w_500_380, w_500_381, w_500_382, w_500_383, w_500_384, w_500_385, w_500_386, w_500_387, w_500_388, w_500_389, w_500_390, w_500_391, w_500_392, w_500_393, w_500_394, w_500_395, w_500_396, w_500_397, w_500_398, w_500_399, w_500_400, w_500_401, w_500_402, w_500_403, w_500_404, w_500_405, w_500_406, w_500_407, w_500_408, w_500_409, w_500_410, w_500_411, w_500_412, w_500_413, w_500_414, w_500_415, w_500_416, w_500_417, w_500_418, w_500_419, w_500_420, w_500_421, w_500_422, w_500_423, w_500_424, w_500_425, w_500_426, w_500_427, w_500_428, w_500_429, w_500_430, w_500_431, w_500_432, w_500_433, w_500_434, w_500_435, w_500_436, w_500_437, w_500_438, w_500_439, w_500_440, w_500_441, w_500_442, w_500_443, w_500_444, w_500_445, w_500_446, w_500_447, w_500_448, w_500_449, w_500_450, w_500_451, w_500_452, w_500_453, w_500_454, w_500_455, w_500_456, w_500_457, w_500_458, w_500_459, w_500_460, w_500_461, w_500_462, w_500_463, w_500_464;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_005);
  nand2 I001_004(w_001_004, w_000_006, w_000_007);
  nand2 I001_005(w_001_005, w_000_008, w_000_009);
  not1 I001_006(w_001_006, w_000_010);
  nand2 I002_000(w_002_000, w_000_011, w_001_002);
  not1 I002_001(w_002_001, w_000_012);
  nand2 I002_002(w_002_002, w_001_002, w_000_013);
  not1 I002_003(w_002_003, w_001_006);
  or2  I002_004(w_002_004, w_000_011, w_000_014);
  or2  I002_005(w_002_005, w_001_006, w_000_015);
  not1 I002_006(w_002_006, w_000_016);
  not1 I002_007(w_002_007, w_001_005);
  nand2 I002_008(w_002_008, w_000_017, w_001_005);
  not1 I002_009(w_002_009, w_000_018);
  or2  I002_010(w_002_010, w_001_000, w_001_003);
  or2  I002_011(w_002_011, w_001_000, w_000_019);
  not1 I002_012(w_002_012, w_001_006);
  nand2 I002_013(w_002_013, w_000_020, w_001_005);
  nand2 I002_014(w_002_014, w_000_021, w_000_022);
  and2 I002_015(w_002_015, w_001_004, w_000_023);
  and2 I002_016(w_002_016, w_000_024, w_000_025);
  and2 I002_017(w_002_017, w_000_026, w_000_027);
  nand2 I002_018(w_002_018, w_000_028, w_000_029);
  or2  I002_019(w_002_019, w_001_003, w_001_002);
  and2 I002_020(w_002_020, w_000_030, w_000_031);
  or2  I002_021(w_002_021, w_001_000, w_000_032);
  and2 I002_022(w_002_022, w_001_003, w_001_006);
  nand2 I002_023(w_002_023, w_001_000, w_001_006);
  or2  I002_024(w_002_024, w_001_002, w_001_005);
  nand2 I002_025(w_002_025, w_001_005, w_000_033);
  and2 I002_026(w_002_026, w_001_003, w_001_004);
  and2 I002_027(w_002_027, w_000_034, w_000_035);
  nand2 I003_000(w_003_000, w_002_021, w_002_003);
  or2  I003_001(w_003_001, w_002_015, w_001_005);
  and2 I003_002(w_003_002, w_001_000, w_002_012);
  and2 I003_003(w_003_003, w_001_004, w_002_019);
  nand2 I003_004(w_003_004, w_002_001, w_000_036);
  and2 I003_005(w_003_005, w_002_017, w_001_002);
  nand2 I003_006(w_003_006, w_000_037, w_002_003);
  or2  I003_007(w_003_007, w_001_004, w_001_003);
  and2 I003_008(w_003_008, w_000_011, w_000_029);
  and2 I003_009(w_003_009, w_001_002, w_001_001);
  not1 I003_010(w_003_010, w_002_004);
  and2 I003_011(w_003_011, w_001_002, w_000_038);
  or2  I003_012(w_003_012, w_002_020, w_002_019);
  not1 I003_013(w_003_013, w_002_014);
  nand2 I003_014(w_003_014, w_001_001, w_001_006);
  or2  I003_015(w_003_015, w_002_006, w_001_001);
  not1 I003_016(w_003_016, w_000_039);
  or2  I003_017(w_003_017, w_000_040, w_001_005);
  nand2 I003_018(w_003_018, w_002_020, w_002_007);
  not1 I003_019(w_003_019, w_002_004);
  not1 I003_020(w_003_020, w_002_002);
  or2  I003_021(w_003_021, w_001_000, w_000_041);
  or2  I003_022(w_003_022, w_000_042, w_001_000);
  not1 I003_023(w_003_023, w_002_012);
  and2 I003_024(w_003_024, w_000_043, w_002_025);
  not1 I003_025(w_003_025, w_002_016);
  and2 I003_026(w_003_026, w_002_007, w_000_044);
  and2 I003_027(w_003_027, w_002_025, w_002_017);
  not1 I003_028(w_003_028, w_001_002);
  and2 I003_029(w_003_029, w_000_045, w_002_007);
  and2 I003_030(w_003_030, w_000_046, w_001_000);
  not1 I003_031(w_003_031, w_001_006);
  not1 I003_032(w_003_032, w_002_004);
  not1 I003_033(w_003_033, w_002_012);
  not1 I003_034(w_003_034, w_000_047);
  or2  I003_035(w_003_035, w_000_048, w_000_049);
  and2 I003_036(w_003_036, w_001_004, w_000_009);
  and2 I003_037(w_003_037, w_002_006, w_002_010);
  or2  I003_038(w_003_038, w_001_001, w_001_003);
  nand2 I003_039(w_003_039, w_001_004, w_002_019);
  nand2 I003_040(w_003_040, w_002_027, w_002_004);
  nand2 I003_041(w_003_041, w_002_008, w_001_000);
  and2 I003_042(w_003_042, w_001_003, w_002_025);
  not1 I003_043(w_003_043, w_002_012);
  and2 I003_044(w_003_044, w_002_014, w_001_000);
  not1 I003_045(w_003_045, w_001_000);
  not1 I003_046(w_003_046, w_002_017);
  not1 I003_047(w_003_047, w_002_024);
  not1 I003_048(w_003_048, w_002_025);
  nand2 I003_049(w_003_049, w_001_001, w_001_004);
  and2 I003_050(w_003_050, w_002_017, w_000_050);
  not1 I003_051(w_003_051, w_001_003);
  not1 I003_052(w_003_052, w_002_020);
  or2  I003_053(w_003_053, w_001_002, w_001_004);
  or2  I003_054(w_003_054, w_001_002, w_000_051);
  and2 I003_055(w_003_055, w_001_006, w_002_004);
  or2  I003_056(w_003_056, w_000_052, w_000_053);
  and2 I003_057(w_003_057, w_000_054, w_000_036);
  and2 I003_058(w_003_058, w_001_003, w_000_055);
  or2  I003_059(w_003_059, w_002_026, w_000_056);
  not1 I003_060(w_003_060, w_002_001);
  and2 I003_061(w_003_061, w_000_057, w_002_025);
  not1 I003_062(w_003_062, w_001_005);
  nand2 I003_063(w_003_063, w_002_001, w_001_004);
  or2  I003_064(w_003_064, w_002_020, w_001_006);
  or2  I003_065(w_003_065, w_000_058, w_000_059);
  or2  I003_066(w_003_066, w_000_060, w_002_027);
  not1 I003_067(w_003_067, w_002_000);
  not1 I003_068(w_003_068, w_002_001);
  nand2 I003_069(w_003_069, w_001_004, w_002_008);
  nand2 I003_070(w_003_070, w_002_013, w_002_010);
  nand2 I003_071(w_003_071, w_002_007, w_002_003);
  and2 I003_072(w_003_072, w_000_061, w_000_062);
  or2  I003_073(w_003_073, w_000_063, w_001_000);
  nand2 I003_074(w_003_074, w_000_064, w_001_002);
  or2  I003_075(w_003_075, w_000_065, w_001_005);
  nand2 I003_076(w_003_076, w_002_004, w_000_066);
  not1 I003_077(w_003_077, w_002_013);
  or2  I003_078(w_003_078, w_002_008, w_002_014);
  and2 I003_079(w_003_079, w_000_023, w_002_025);
  or2  I003_080(w_003_080, w_000_067, w_002_003);
  or2  I003_081(w_003_081, w_000_068, w_001_003);
  or2  I003_082(w_003_082, w_002_000, w_000_069);
  and2 I003_083(w_003_083, w_001_002, w_000_070);
  not1 I003_084(w_003_084, w_001_003);
  not1 I003_085(w_003_085, w_001_005);
  not1 I003_086(w_003_086, w_002_022);
  nand2 I003_087(w_003_087, w_000_071, w_001_000);
  nand2 I003_088(w_003_088, w_002_022, w_000_072);
  and2 I003_089(w_003_089, w_002_020, w_000_073);
  or2  I003_090(w_003_090, w_000_074, w_002_001);
  and2 I003_091(w_003_091, w_000_075, w_001_002);
  not1 I003_092(w_003_092, w_001_004);
  and2 I003_093(w_003_093, w_000_076, w_001_006);
  or2  I003_094(w_003_094, w_000_059, w_002_018);
  or2  I003_095(w_003_095, w_000_077, w_002_009);
  or2  I003_096(w_003_096, w_000_078, w_001_002);
  or2  I003_097(w_003_097, w_001_002, w_000_079);
  nand2 I003_098(w_003_098, w_002_018, w_002_024);
  not1 I003_099(w_003_099, w_002_017);
  or2  I003_100(w_003_100, w_000_080, w_001_003);
  or2  I003_101(w_003_101, w_001_006, w_001_003);
  or2  I004_000(w_004_000, w_003_023, w_002_014);
  not1 I004_001(w_004_001, w_000_081);
  or2  I004_002(w_004_002, w_003_021, w_001_004);
  nand2 I004_003(w_004_003, w_003_043, w_003_021);
  or2  I004_004(w_004_004, w_000_054, w_002_014);
  or2  I004_005(w_004_005, w_001_002, w_000_002);
  nand2 I004_006(w_004_006, w_003_092, w_000_082);
  and2 I004_007(w_004_007, w_002_021, w_002_026);
  and2 I004_008(w_004_008, w_003_069, w_001_001);
  and2 I004_009(w_004_009, w_000_083, w_003_055);
  or2  I004_010(w_004_010, w_000_084, w_003_025);
  not1 I004_011(w_004_011, w_000_060);
  not1 I004_012(w_004_012, w_001_000);
  nand2 I004_014(w_004_014, w_003_047, w_002_005);
  and2 I004_015(w_004_015, w_001_005, w_001_004);
  not1 I004_016(w_004_016, w_002_021);
  not1 I004_017(w_004_017, w_001_004);
  not1 I004_018(w_004_018, w_001_003);
  or2  I004_019(w_004_019, w_003_074, w_002_017);
  nand2 I004_020(w_004_020, w_001_003, w_003_088);
  nand2 I004_021(w_004_021, w_002_008, w_002_017);
  not1 I004_022(w_004_022, w_003_035);
  nand2 I004_023(w_004_023, w_001_002, w_001_006);
  or2  I004_024(w_004_024, w_003_006, w_002_021);
  and2 I004_025(w_004_025, w_003_055, w_002_022);
  not1 I004_026(w_004_026, w_000_071);
  or2  I004_027(w_004_027, w_001_003, w_000_086);
  or2  I004_028(w_004_028, w_002_004, w_003_077);
  not1 I004_029(w_004_029, w_003_037);
  or2  I004_030(w_004_030, w_000_087, w_002_011);
  or2  I004_031(w_004_031, w_000_088, w_001_004);
  and2 I004_032(w_004_032, w_003_066, w_002_015);
  nand2 I004_034(w_004_034, w_001_004, w_000_090);
  not1 I004_036(w_004_036, w_002_007);
  nand2 I004_037(w_004_037, w_002_002, w_001_004);
  nand2 I004_038(w_004_038, w_002_019, w_000_082);
  nand2 I004_039(w_004_039, w_000_091, w_002_023);
  and2 I004_043(w_004_043, w_003_018, w_000_092);
  not1 I004_044(w_004_044, w_003_015);
  or2  I004_046(w_004_046, w_002_005, w_003_051);
  or2  I004_047(w_004_047, w_003_051, w_000_093);
  or2  I004_048(w_004_048, w_000_084, w_000_094);
  not1 I004_050(w_004_050, w_003_052);
  nand2 I004_051(w_004_051, w_001_003, w_002_010);
  and2 I004_052(w_004_052, w_000_095, w_003_000);
  not1 I004_053(w_004_053, w_001_004);
  or2  I004_054(w_004_054, w_002_002, w_001_006);
  nand2 I004_057(w_004_057, w_002_002, w_002_019);
  or2  I004_058(w_004_058, w_001_004, w_003_016);
  or2  I004_059(w_004_059, w_002_013, w_003_007);
  and2 I004_060(w_004_060, w_001_005, w_002_000);
  nand2 I004_061(w_004_061, w_001_004, w_002_013);
  not1 I004_062(w_004_062, w_003_057);
  nand2 I004_065(w_004_065, w_000_097, w_001_000);
  nand2 I004_066(w_004_066, w_000_098, w_003_083);
  not1 I004_067(w_004_067, w_001_003);
  and2 I004_069(w_004_069, w_000_099, w_000_025);
  and2 I004_070(w_004_070, w_003_025, w_002_024);
  and2 I004_071(w_004_071, w_002_003, w_001_001);
  not1 I004_072(w_004_072, w_001_002);
  nand2 I004_076(w_004_076, w_002_017, w_003_049);
  and2 I004_078(w_004_078, w_002_001, w_001_005);
  or2  I004_080(w_004_080, w_003_055, w_002_004);
  or2  I004_081(w_004_081, w_001_004, w_000_101);
  and2 I004_082(w_004_082, w_003_072, w_001_000);
  and2 I004_083(w_004_083, w_002_000, w_000_093);
  not1 I004_084(w_004_084, w_001_006);
  and2 I004_085(w_004_085, w_002_025, w_000_102);
  or2  I004_086(w_004_086, w_003_004, w_003_076);
  or2  I004_087(w_004_087, w_001_005, w_003_028);
  or2  I004_088(w_004_088, w_003_077, w_001_004);
  or2  I004_089(w_004_089, w_002_024, w_001_006);
  or2  I004_091(w_004_091, w_002_005, w_003_006);
  nand2 I004_094(w_004_094, w_000_104, w_000_090);
  or2  I004_095(w_004_095, w_002_016, w_001_004);
  or2  I004_096(w_004_096, w_001_004, w_003_045);
  and2 I004_097(w_004_097, w_000_006, w_002_027);
  and2 I004_098(w_004_098, w_001_004, w_002_020);
  or2  I004_100(w_004_100, w_000_105, w_000_106);
  nand2 I004_102(w_004_102, w_003_061, w_003_050);
  or2  I004_103(w_004_103, w_001_003, w_001_004);
  nand2 I004_104(w_004_104, w_001_005, w_003_048);
  nand2 I004_105(w_004_105, w_001_005, w_001_002);
  or2  I004_106(w_004_106, w_003_053, w_001_006);
  and2 I004_107(w_004_107, w_000_107, w_003_082);
  or2  I004_109(w_004_109, w_001_000, w_003_050);
  and2 I004_110(w_004_110, w_002_019, w_000_042);
  and2 I004_111(w_004_111, w_003_011, w_001_001);
  or2  I004_112(w_004_112, w_002_023, w_000_109);
  nand2 I004_113(w_004_113, w_001_000, w_000_110);
  or2  I004_114(w_004_114, w_003_064, w_003_059);
  and2 I004_115(w_004_115, w_000_111, w_002_004);
  and2 I004_117(w_004_117, w_003_071, w_003_064);
  or2  I004_118(w_004_118, w_001_006, w_002_001);
  or2  I004_120(w_004_120, w_000_113, w_002_001);
  nand2 I004_121(w_004_121, w_002_020, w_002_004);
  nand2 I004_122(w_004_122, w_000_114, w_002_010);
  and2 I004_124(w_004_124, w_003_030, w_001_003);
  nand2 I004_125(w_004_125, w_002_024, w_001_001);
  nand2 I004_127(w_004_127, w_001_003, w_000_115);
  nand2 I004_128(w_004_128, w_003_024, w_000_116);
  or2  I004_130(w_004_130, w_002_009, w_002_013);
  nand2 I004_131(w_004_131, w_003_075, w_002_009);
  nand2 I004_132(w_004_132, w_003_033, w_000_117);
  not1 I004_133(w_004_133, w_002_015);
  or2  I004_134(w_004_134, w_003_084, w_001_004);
  not1 I004_135(w_004_135, w_001_002);
  not1 I004_136(w_004_136, w_003_069);
  nand2 I004_137(w_004_137, w_003_038, w_002_020);
  and2 I004_138(w_004_138, w_003_055, w_003_010);
  or2  I004_139(w_004_139, w_000_118, w_001_005);
  nand2 I004_141(w_004_141, w_003_047, w_001_002);
  nand2 I004_142(w_004_142, w_002_001, w_002_005);
  not1 I004_143(w_004_143, w_001_005);
  and2 I004_144(w_004_144, w_003_057, w_001_004);
  nand2 I004_147(w_004_147, w_000_045, w_002_007);
  nand2 I004_148(w_004_148, w_003_089, w_002_017);
  not1 I004_149(w_004_149, w_000_121);
  not1 I004_152(w_004_152, w_002_011);
  nand2 I004_154(w_004_154, w_001_006, w_001_002);
  and2 I004_155(w_004_155, w_001_000, w_003_014);
  nand2 I004_156(w_004_156, w_003_069, w_003_097);
  and2 I004_157(w_004_157, w_000_071, w_000_124);
  not1 I004_159(w_004_159, w_002_004);
  not1 I004_160(w_004_160, w_000_124);
  or2  I004_161(w_004_161, w_001_004, w_003_064);
  or2  I004_163(w_004_163, w_002_027, w_001_004);
  not1 I004_164(w_004_164, w_002_019);
  and2 I004_166(w_004_166, w_001_003, w_003_040);
  nand2 I004_167(w_004_167, w_002_001, w_003_040);
  or2  I004_168(w_004_168, w_000_125, w_002_018);
  and2 I004_172(w_004_172, w_003_072, w_000_096);
  not1 I004_173(w_004_173, w_003_090);
  and2 I004_175(w_004_175, w_000_128, w_003_082);
  and2 I004_178(w_004_178, w_001_006, w_000_129);
  or2  I004_179(w_004_179, w_000_130, w_003_059);
  nand2 I004_180(w_004_180, w_000_131, w_002_024);
  nand2 I004_181(w_004_181, w_003_043, w_003_030);
  nand2 I004_182(w_004_182, w_000_132, w_002_022);
  or2  I004_183(w_004_183, w_003_091, w_003_101);
  and2 I004_184(w_004_184, w_003_061, w_003_023);
  nand2 I004_186(w_004_186, w_001_004, w_000_134);
  nand2 I004_187(w_004_187, w_003_030, w_000_135);
  and2 I004_188(w_004_188, w_000_098, w_002_018);
  and2 I004_189(w_004_189, w_003_098, w_003_010);
  or2  I004_190(w_004_190, w_003_040, w_002_014);
  or2  I004_191(w_004_191, w_000_136, w_001_004);
  or2  I004_192(w_004_192, w_000_047, w_000_016);
  not1 I004_193(w_004_193, w_000_137);
  or2  I004_194(w_004_194, w_000_053, w_001_005);
  nand2 I004_195(w_004_195, w_003_043, w_003_090);
  nand2 I004_198(w_004_198, w_001_003, w_000_139);
  not1 I004_199(w_004_199, w_001_005);
  or2  I004_201(w_004_201, w_003_032, w_000_140);
  or2  I004_202(w_004_202, w_003_061, w_002_010);
  not1 I004_203(w_004_203, w_000_116);
  or2  I004_204(w_004_204, w_001_000, w_001_002);
  nand2 I004_206(w_004_206, w_001_005, w_000_062);
  not1 I004_209(w_004_209, w_000_040);
  and2 I004_210(w_004_210, w_002_018, w_001_000);
  nand2 I004_211(w_004_211, w_002_018, w_000_144);
  not1 I004_213(w_004_213, w_000_034);
  nand2 I004_214(w_004_214, w_002_026, w_001_005);
  nand2 I004_215(w_004_215, w_000_145, w_000_146);
  or2  I004_216(w_004_216, w_003_012, w_001_000);
  or2  I004_217(w_004_217, w_003_055, w_002_005);
  or2  I004_219(w_004_219, w_000_128, w_003_004);
  and2 I004_221(w_004_221, w_003_058, w_003_000);
  nand2 I004_222(w_004_222, w_003_030, w_000_149);
  not1 I004_223(w_004_223, w_001_000);
  nand2 I004_224(w_004_224, w_000_150, w_001_003);
  not1 I004_225(w_004_225, w_002_024);
  nand2 I004_226(w_004_226, w_003_034, w_003_043);
  or2  I004_227(w_004_227, w_003_057, w_000_151);
  or2  I004_228(w_004_228, w_003_091, w_001_000);
  not1 I004_230(w_004_230, w_003_072);
  or2  I004_232(w_004_232, w_000_154, w_003_077);
  and2 I004_233(w_004_233, w_002_007, w_003_010);
  and2 I004_234(w_004_234, w_002_019, w_000_067);
  or2  I004_237(w_004_237, w_003_088, w_000_147);
  or2  I004_238(w_004_238, w_001_006, w_002_000);
  and2 I004_239(w_004_239, w_003_051, w_003_062);
  or2  I004_240(w_004_240, w_000_153, w_000_052);
  and2 I004_241(w_004_241, w_001_001, w_003_075);
  nand2 I004_243(w_004_243, w_002_004, w_001_002);
  nand2 I004_244(w_004_244, w_002_020, w_003_017);
  and2 I004_245(w_004_245, w_003_014, w_003_019);
  not1 I004_246(w_004_246, w_000_011);
  nand2 I004_247(w_004_247, w_001_000, w_000_156);
  and2 I004_249(w_004_249, w_001_005, w_003_081);
  not1 I004_250(w_004_250, w_001_001);
  or2  I004_251(w_004_251, w_003_021, w_000_044);
  not1 I004_252(w_004_252, w_000_012);
  or2  I004_253(w_004_253, w_003_043, w_002_002);
  not1 I004_254(w_004_254, w_003_077);
  not1 I004_255(w_004_255, w_001_002);
  not1 I004_256(w_004_256, w_003_005);
  not1 I004_257(w_004_257, w_003_014);
  nand2 I004_259(w_004_259, w_003_001, w_000_158);
  and2 I004_260(w_004_260, w_002_004, w_000_004);
  not1 I004_263(w_004_263, w_002_025);
  or2  I004_265(w_004_265, w_003_094, w_000_159);
  not1 I004_267(w_004_267, w_000_131);
  or2  I004_268(w_004_268, w_000_160, w_002_010);
  not1 I004_269(w_004_269, w_001_003);
  not1 I004_271(w_004_271, w_000_161);
  nand2 I004_272(w_004_272, w_001_000, w_002_009);
  and2 I004_273(w_004_273, w_000_162, w_001_006);
  or2  I004_274(w_004_274, w_001_006, w_002_016);
  nand2 I004_275(w_004_275, w_002_022, w_001_000);
  and2 I004_276(w_004_276, w_002_002, w_001_004);
  nand2 I004_277(w_004_277, w_000_050, w_001_002);
  and2 I004_278(w_004_278, w_000_163, w_000_134);
  nand2 I004_279(w_004_279, w_001_000, w_001_005);
  not1 I004_280(w_004_280, w_002_023);
  not1 I004_282(w_004_282, w_000_165);
  not1 I004_283(w_004_283, w_002_017);
  not1 I004_285(w_004_285, w_001_004);
  not1 I004_286(w_004_286, w_003_017);
  or2  I004_287(w_004_287, w_003_000, w_000_048);
  nand2 I004_289(w_004_289, w_000_166, w_001_000);
  and2 I004_290(w_004_290, w_000_167, w_002_001);
  and2 I004_291(w_004_291, w_000_168, w_001_003);
  nand2 I004_292(w_004_292, w_002_005, w_002_002);
  not1 I004_293(w_004_293, w_003_063);
  nand2 I004_295(w_004_295, w_000_170, w_002_012);
  not1 I004_296(w_004_296, w_000_171);
  not1 I004_297(w_004_297, w_000_023);
  and2 I004_300(w_004_300, w_001_001, w_003_050);
  or2  I004_301(w_004_301, w_002_011, w_001_004);
  not1 I004_302(w_004_302, w_002_013);
  or2  I004_303(w_004_303, w_002_000, w_001_000);
  not1 I004_304(w_004_304, w_001_001);
  nand2 I004_305(w_004_305, w_002_023, w_001_001);
  not1 I004_307(w_004_307, w_000_172);
  or2  I004_308(w_004_308, w_002_024, w_003_091);
  or2  I004_309(w_004_309, w_002_023, w_003_008);
  and2 I004_310(w_004_310, w_002_012, w_001_004);
  not1 I004_311(w_004_311, w_002_019);
  not1 I004_312(w_004_312, w_000_130);
  nand2 I004_313(w_004_313, w_001_004, w_002_027);
  or2  I004_314(w_004_314, w_000_173, w_001_001);
  nand2 I004_315(w_004_315, w_003_023, w_003_078);
  and2 I004_316(w_004_316, w_001_001, w_000_174);
  and2 I004_317(w_004_317, w_002_009, w_002_013);
  and2 I004_318(w_004_318, w_000_052, w_002_013);
  not1 I004_319(w_004_319, w_001_002);
  or2  I004_320(w_004_320, w_003_041, w_002_011);
  nand2 I004_321(w_004_321, w_000_175, w_003_039);
  or2  I004_322(w_004_322, w_002_016, w_001_005);
  and2 I004_323(w_004_323, w_001_006, w_000_063);
  not1 I004_324(w_004_324, w_002_008);
  not1 I004_325(w_004_325, w_003_036);
  and2 I004_327(w_004_327, w_000_039, w_002_027);
  nand2 I004_328(w_004_328, w_002_001, w_002_026);
  not1 I004_329(w_004_329, w_000_176);
  and2 I004_330(w_004_330, w_003_054, w_001_003);
  not1 I004_331(w_004_331, w_001_001);
  or2  I004_332(w_004_332, w_001_005, w_000_142);
  not1 I004_333(w_004_333, w_000_065);
  not1 I004_336(w_004_336, w_000_178);
  not1 I004_338(w_004_338, w_000_179);
  not1 I004_339(w_004_339, w_002_026);
  or2  I004_340(w_004_340, w_003_057, w_003_087);
  or2  I004_341(w_004_341, w_001_005, w_002_008);
  or2  I004_342(w_004_342, w_003_086, w_003_035);
  and2 I004_343(w_004_343, w_003_047, w_001_001);
  or2  I004_344(w_004_344, w_000_096, w_003_050);
  not1 I004_345(w_004_345, w_003_039);
  or2  I004_346(w_004_346, w_001_006, w_002_025);
  not1 I004_347(w_004_347, w_001_005);
  and2 I004_348(w_004_348, w_002_008, w_002_015);
  or2  I004_349(w_004_349, w_002_019, w_000_180);
  nand2 I004_350(w_004_350, w_000_181, w_000_182);
  nand2 I004_351(w_004_351, w_001_005, w_002_009);
  or2  I004_352(w_004_352, w_001_002, w_002_026);
  or2  I004_353(w_004_353, w_000_047, w_003_020);
  and2 I004_354(w_004_354, w_003_054, w_000_183);
  or2  I004_356(w_004_356, w_002_002, w_003_057);
  and2 I004_357(w_004_357, w_002_016, w_001_004);
  or2  I004_358(w_004_358, w_003_101, w_003_042);
  not1 I004_359(w_004_359, w_003_087);
  and2 I004_360(w_004_360, w_003_039, w_000_184);
  or2  I004_361(w_004_361, w_000_185, w_001_004);
  not1 I004_362(w_004_362, w_002_001);
  and2 I004_363(w_004_363, w_001_003, w_000_043);
  and2 I004_365(w_004_365, w_000_186, w_003_034);
  not1 I004_366(w_004_366, w_002_008);
  not1 I004_367(w_004_367, w_001_004);
  not1 I004_368(w_004_368, w_000_056);
  not1 I004_369(w_004_369, w_001_000);
  or2  I004_370(w_004_370, w_003_071, w_003_074);
  and2 I004_371(w_004_371, w_003_090, w_003_042);
  nand2 I004_372(w_004_372, w_002_005, w_002_006);
  not1 I004_373(w_004_373, w_002_005);
  not1 I004_374(w_004_374, w_000_008);
  or2  I004_376(w_004_376, w_000_187, w_001_006);
  nand2 I004_378(w_004_378, w_002_025, w_003_007);
  and2 I004_380(w_004_380, w_000_126, w_002_002);
  or2  I004_381(w_004_381, w_002_026, w_003_100);
  and2 I004_383(w_004_383, w_000_069, w_000_188);
  not1 I004_384(w_004_384, w_000_189);
  and2 I004_385(w_004_385, w_003_082, w_000_190);
  nand2 I004_386(w_004_386, w_003_014, w_003_015);
  or2  I004_387(w_004_387, w_002_025, w_002_024);
  nand2 I004_388(w_004_388, w_001_003, w_003_090);
  not1 I004_389(w_004_389, w_000_057);
  or2  I004_393(w_004_393, w_002_001, w_003_027);
  and2 I004_394(w_004_394, w_002_024, w_003_055);
  not1 I004_395(w_004_395, w_001_005);
  nand2 I004_396(w_004_396, w_000_191, w_000_055);
  or2  I004_397(w_004_397, w_002_020, w_002_008);
  or2  I004_398(w_004_398, w_000_050, w_001_000);
  or2  I004_399(w_004_399, w_002_017, w_002_004);
  not1 I004_400(w_004_400, w_002_025);
  not1 I004_401(w_004_401, w_000_054);
  or2  I004_402(w_004_402, w_003_012, w_002_008);
  nand2 I004_405(w_004_405, w_001_006, w_000_186);
  or2  I004_406(w_004_406, w_003_075, w_003_071);
  or2  I004_407(w_004_407, w_001_005, w_003_047);
  nand2 I004_408(w_004_408, w_000_024, w_003_091);
  and2 I004_410(w_004_410, w_002_020, w_003_096);
  nand2 I004_412(w_004_412, w_002_006, w_002_002);
  or2  I004_413(w_004_413, w_003_075, w_002_026);
  not1 I004_415(w_004_415, w_002_012);
  and2 I004_416(w_004_416, w_001_006, w_000_035);
  not1 I004_417(w_004_417, w_003_029);
  and2 I004_418(w_004_418, w_002_013, w_001_003);
  and2 I004_419(w_004_419, w_000_192, w_003_002);
  not1 I004_421(w_004_421, w_000_156);
  not1 I004_424(w_004_424, w_002_002);
  not1 I004_425(w_004_425, w_002_022);
  and2 I004_426(w_004_426, w_003_080, w_001_002);
  and2 I004_427(w_004_427, w_000_193, w_002_020);
  or2  I004_428(w_004_428, w_003_041, w_002_014);
  and2 I004_429(w_004_429, w_002_006, w_001_005);
  and2 I004_430(w_004_430, w_003_080, w_003_095);
  and2 I004_431(w_004_431, w_001_006, w_002_011);
  and2 I004_432(w_004_432, w_002_014, w_000_043);
  not1 I004_433(w_004_433, w_000_194);
  nand2 I004_435(w_004_435, w_003_011, w_003_017);
  or2  I004_436(w_004_436, w_001_006, w_001_005);
  and2 I004_438(w_004_438, w_002_021, w_000_029);
  and2 I004_439(w_004_439, w_000_196, w_002_000);
  and2 I004_440(w_004_440, w_002_006, w_000_197);
  and2 I004_441(w_004_441, w_003_063, w_003_017);
  or2  I004_442(w_004_442, w_001_005, w_002_018);
  or2  I004_444(w_004_444, w_003_046, w_002_012);
  or2  I004_445(w_004_445, w_002_012, w_002_008);
  or2  I004_446(w_004_446, w_002_023, w_003_062);
  nand2 I004_447(w_004_447, w_003_061, w_002_003);
  and2 I004_448(w_004_448, w_003_064, w_000_026);
  not1 I004_449(w_004_449, w_000_198);
  not1 I004_451(w_004_451, w_001_000);
  and2 I004_452(w_004_452, w_003_059, w_002_004);
  not1 I004_454(w_004_454, w_003_051);
  and2 I004_455(w_004_455, w_002_016, w_000_200);
  and2 I004_456(w_004_456, w_002_017, w_001_006);
  not1 I004_457(w_004_457, w_000_201);
  or2  I004_458(w_004_458, w_003_100, w_002_026);
  not1 I004_459(w_004_459, w_001_003);
  and2 I004_460(w_004_460, w_001_006, w_000_202);
  not1 I004_462(w_004_462, w_002_015);
  and2 I004_463(w_004_463, w_002_011, w_003_028);
  or2  I004_464(w_004_464, w_000_135, w_003_046);
  and2 I004_465(w_004_465, w_003_055, w_003_037);
  and2 I004_467(w_004_467, w_000_203, w_001_003);
  or2  I004_468(w_004_468, w_003_099, w_003_017);
  not1 I004_469(w_004_469, w_003_071);
  or2  I004_470(w_004_470, w_002_014, w_002_006);
  or2  I004_471(w_004_471, w_001_004, w_000_117);
  not1 I004_472(w_004_472, w_002_011);
  not1 I004_473(w_004_473, w_001_000);
  not1 I004_474(w_004_474, w_001_001);
  not1 I005_000(w_005_000, w_000_204);
  not1 I005_001(w_005_001, w_002_020);
  and2 I005_002(w_005_002, w_003_084, w_004_023);
  not1 I005_003(w_005_003, w_000_205);
  nand2 I005_004(w_005_004, w_001_002, w_002_010);
  nand2 I005_005(w_005_005, w_004_352, w_004_393);
  not1 I005_006(w_005_006, w_002_004);
  or2  I005_007(w_005_007, w_004_413, w_002_022);
  and2 I005_008(w_005_008, w_002_004, w_001_004);
  or2  I005_009(w_005_009, w_001_003, w_002_022);
  not1 I005_010(w_005_010, w_004_296);
  or2  I005_011(w_005_011, w_000_206, w_001_005);
  not1 I005_012(w_005_012, w_002_004);
  and2 I005_013(w_005_013, w_002_007, w_001_000);
  and2 I005_014(w_005_014, w_000_207, w_002_025);
  nand2 I005_015(w_005_015, w_000_057, w_004_048);
  not1 I005_016(w_005_016, w_001_001);
  or2  I005_017(w_005_017, w_003_054, w_002_021);
  nand2 I005_018(w_005_018, w_004_324, w_002_002);
  not1 I005_019(w_005_019, w_004_139);
  not1 I005_020(w_005_020, w_004_342);
  or2  I005_021(w_005_021, w_002_010, w_002_008);
  not1 I005_022(w_005_022, w_000_075);
  not1 I005_023(w_005_023, w_000_160);
  not1 I005_024(w_005_024, w_000_123);
  not1 I005_025(w_005_025, w_000_208);
  and2 I005_026(w_005_026, w_004_149, w_002_025);
  or2  I005_027(w_005_027, w_004_448, w_001_003);
  nand2 I005_028(w_005_028, w_002_012, w_004_459);
  not1 I005_029(w_005_029, w_003_082);
  not1 I005_030(w_005_030, w_002_027);
  not1 I005_031(w_005_031, w_001_001);
  not1 I005_032(w_005_032, w_000_109);
  or2  I005_033(w_005_033, w_000_209, w_002_005);
  not1 I005_034(w_005_034, w_003_085);
  and2 I005_035(w_005_035, w_003_033, w_004_011);
  and2 I005_036(w_005_036, w_003_062, w_001_005);
  nand2 I005_037(w_005_037, w_000_210, w_001_002);
  and2 I005_038(w_005_038, w_003_071, w_002_014);
  or2  I005_039(w_005_039, w_000_211, w_003_094);
  nand2 I005_040(w_005_040, w_002_017, w_004_393);
  and2 I005_041(w_005_041, w_000_212, w_003_096);
  and2 I005_042(w_005_042, w_002_011, w_004_026);
  or2  I005_043(w_005_043, w_001_002, w_003_062);
  or2  I005_044(w_005_044, w_001_006, w_001_003);
  nand2 I005_045(w_005_045, w_004_280, w_002_002);
  nand2 I005_046(w_005_046, w_003_057, w_001_005);
  or2  I005_047(w_005_047, w_003_066, w_001_000);
  or2  I005_048(w_005_048, w_002_010, w_000_213);
  and2 I005_049(w_005_049, w_003_029, w_004_124);
  nand2 I005_050(w_005_050, w_003_037, w_000_214);
  nand2 I005_052(w_005_052, w_000_155, w_002_016);
  nand2 I005_053(w_005_053, w_001_000, w_003_036);
  and2 I005_055(w_005_055, w_000_072, w_002_003);
  and2 I005_056(w_005_056, w_002_026, w_004_098);
  and2 I005_057(w_005_057, w_002_005, w_003_098);
  nand2 I005_058(w_005_058, w_002_014, w_000_114);
  nand2 I005_059(w_005_059, w_001_003, w_000_215);
  and2 I005_060(w_005_060, w_003_075, w_000_216);
  not1 I005_061(w_005_061, w_002_016);
  nand2 I005_062(w_005_062, w_000_217, w_000_218);
  not1 I005_064(w_005_064, w_003_002);
  nand2 I005_065(w_005_065, w_003_044, w_000_219);
  or2  I005_066(w_005_066, w_001_006, w_001_005);
  nand2 I005_067(w_005_067, w_003_031, w_003_017);
  and2 I005_068(w_005_068, w_002_022, w_001_001);
  or2  I005_069(w_005_069, w_001_003, w_000_190);
  and2 I005_070(w_005_070, w_002_024, w_003_057);
  not1 I005_071(w_005_071, w_001_001);
  and2 I005_072(w_005_072, w_003_040, w_002_001);
  nand2 I005_073(w_005_073, w_001_004, w_003_023);
  and2 I005_074(w_005_074, w_003_050, w_003_010);
  not1 I005_075(w_005_075, w_004_470);
  nand2 I005_076(w_005_076, w_000_220, w_000_040);
  and2 I005_077(w_005_077, w_004_280, w_003_025);
  nand2 I005_078(w_005_078, w_004_004, w_003_019);
  or2  I005_080(w_005_080, w_004_083, w_002_000);
  nand2 I005_081(w_005_081, w_000_196, w_000_054);
  not1 I005_082(w_005_082, w_004_256);
  not1 I005_083(w_005_083, w_004_296);
  not1 I005_084(w_005_084, w_000_221);
  and2 I005_085(w_005_085, w_002_016, w_002_022);
  nand2 I005_086(w_005_086, w_003_033, w_003_084);
  nand2 I005_087(w_005_087, w_002_000, w_000_222);
  not1 I005_088(w_005_088, w_000_223);
  or2  I005_089(w_005_089, w_001_004, w_003_093);
  and2 I005_090(w_005_090, w_004_389, w_003_027);
  nand2 I005_091(w_005_091, w_003_048, w_000_224);
  and2 I005_092(w_005_092, w_004_130, w_001_003);
  nand2 I005_093(w_005_093, w_001_004, w_000_225);
  not1 I005_094(w_005_094, w_002_008);
  and2 I005_095(w_005_095, w_002_013, w_002_018);
  and2 I005_096(w_005_096, w_002_001, w_001_004);
  not1 I005_097(w_005_097, w_001_003);
  or2  I005_098(w_005_098, w_001_000, w_004_069);
  and2 I005_099(w_005_099, w_000_051, w_003_026);
  nand2 I005_100(w_005_100, w_004_072, w_000_226);
  nand2 I005_101(w_005_101, w_004_009, w_004_016);
  not1 I005_103(w_005_103, w_000_227);
  and2 I005_104(w_005_104, w_001_006, w_001_003);
  nand2 I005_105(w_005_105, w_000_228, w_000_167);
  nand2 I005_106(w_005_106, w_003_091, w_002_000);
  or2  I005_107(w_005_107, w_004_107, w_001_004);
  nand2 I005_108(w_005_108, w_003_085, w_003_011);
  not1 I005_109(w_005_109, w_002_010);
  and2 I005_110(w_005_110, w_004_387, w_000_072);
  nand2 I005_111(w_005_111, w_001_005, w_003_038);
  not1 I005_112(w_005_112, w_003_001);
  or2  I005_113(w_005_113, w_002_026, w_003_008);
  nand2 I005_114(w_005_114, w_002_001, w_001_006);
  or2  I005_115(w_005_115, w_004_406, w_003_033);
  nand2 I005_117(w_005_117, w_003_047, w_000_229);
  or2  I005_118(w_005_118, w_003_053, w_001_002);
  and2 I005_119(w_005_119, w_002_022, w_001_005);
  and2 I005_120(w_005_120, w_000_230, w_003_001);
  nand2 I005_121(w_005_121, w_003_069, w_002_004);
  not1 I005_122(w_005_122, w_002_017);
  not1 I005_123(w_005_123, w_000_104);
  or2  I005_124(w_005_124, w_000_207, w_000_231);
  or2  I005_125(w_005_125, w_004_105, w_003_051);
  or2  I005_126(w_005_126, w_001_004, w_004_276);
  nand2 I005_127(w_005_127, w_002_007, w_004_130);
  and2 I005_130(w_005_130, w_000_181, w_003_090);
  and2 I005_132(w_005_132, w_004_023, w_000_232);
  not1 I005_133(w_005_133, w_001_006);
  or2  I005_134(w_005_134, w_003_093, w_001_006);
  or2  I005_135(w_005_135, w_001_002, w_004_180);
  nand2 I005_136(w_005_136, w_004_257, w_001_000);
  not1 I005_137(w_005_137, w_001_003);
  nand2 I005_138(w_005_138, w_002_025, w_000_224);
  not1 I005_139(w_005_139, w_002_023);
  not1 I005_141(w_005_141, w_001_001);
  and2 I005_142(w_005_142, w_002_012, w_001_004);
  or2  I005_143(w_005_143, w_001_000, w_003_099);
  or2  I005_144(w_005_144, w_001_000, w_001_004);
  nand2 I005_145(w_005_145, w_000_026, w_003_024);
  and2 I005_146(w_005_146, w_000_233, w_003_068);
  nand2 I005_147(w_005_147, w_003_076, w_001_001);
  not1 I005_148(w_005_148, w_001_001);
  not1 I005_149(w_005_149, w_000_234);
  and2 I005_150(w_005_150, w_003_060, w_001_004);
  and2 I005_151(w_005_151, w_003_018, w_000_140);
  nand2 I005_152(w_005_152, w_002_018, w_000_222);
  nand2 I005_153(w_005_153, w_000_004, w_003_042);
  nand2 I005_154(w_005_154, w_001_000, w_003_081);
  and2 I005_155(w_005_155, w_002_006, w_001_004);
  nand2 I005_156(w_005_156, w_002_010, w_001_005);
  not1 I005_157(w_005_157, w_000_235);
  not1 I005_158(w_005_158, w_002_002);
  not1 I005_159(w_005_159, w_004_469);
  not1 I005_160(w_005_160, w_004_012);
  and2 I005_161(w_005_161, w_003_041, w_003_051);
  or2  I005_162(w_005_162, w_003_061, w_001_005);
  or2  I005_163(w_005_163, w_001_002, w_004_354);
  not1 I005_164(w_005_164, w_002_024);
  not1 I005_165(w_005_165, w_000_236);
  and2 I005_166(w_005_166, w_001_002, w_001_005);
  or2  I005_167(w_005_167, w_000_189, w_003_100);
  or2  I005_168(w_005_168, w_003_049, w_002_016);
  and2 I005_169(w_005_169, w_000_237, w_001_002);
  or2  I005_170(w_005_170, w_002_003, w_002_026);
  not1 I005_171(w_005_171, w_001_005);
  and2 I005_172(w_005_172, w_004_289, w_004_210);
  or2  I005_173(w_005_173, w_000_001, w_000_238);
  and2 I005_175(w_005_175, w_003_005, w_001_000);
  nand2 I005_176(w_005_176, w_004_471, w_002_007);
  and2 I005_177(w_005_177, w_001_003, w_002_003);
  and2 I005_178(w_005_178, w_000_162, w_002_026);
  nand2 I005_179(w_005_179, w_004_396, w_004_296);
  or2  I005_180(w_005_180, w_004_096, w_002_021);
  nand2 I005_181(w_005_181, w_001_005, w_003_061);
  or2  I005_182(w_005_182, w_002_022, w_002_018);
  not1 I005_184(w_005_184, w_001_003);
  and2 I005_185(w_005_185, w_004_400, w_000_038);
  or2  I005_186(w_005_186, w_000_239, w_001_001);
  not1 I005_187(w_005_187, w_000_216);
  not1 I005_188(w_005_188, w_001_003);
  and2 I005_189(w_005_189, w_004_351, w_004_452);
  and2 I005_190(w_005_190, w_001_003, w_003_058);
  not1 I005_191(w_005_191, w_004_130);
  not1 I005_192(w_005_192, w_002_010);
  nand2 I005_193(w_005_193, w_002_001, w_000_221);
  or2  I005_194(w_005_194, w_000_120, w_001_001);
  not1 I005_195(w_005_195, w_002_004);
  or2  I005_196(w_005_196, w_004_269, w_000_240);
  nand2 I005_197(w_005_197, w_002_024, w_004_309);
  not1 I005_198(w_005_198, w_003_091);
  and2 I005_199(w_005_199, w_000_038, w_002_012);
  or2  I005_200(w_005_200, w_001_006, w_001_002);
  not1 I005_201(w_005_201, w_002_009);
  nand2 I005_203(w_005_203, w_001_001, w_003_088);
  nand2 I005_206(w_005_206, w_001_006, w_000_012);
  and2 I005_207(w_005_207, w_003_058, w_004_038);
  and2 I005_208(w_005_208, w_003_042, w_000_241);
  or2  I005_210(w_005_210, w_002_013, w_000_023);
  nand2 I005_211(w_005_211, w_000_242, w_001_006);
  or2  I005_212(w_005_212, w_000_243, w_002_023);
  not1 I005_213(w_005_213, w_000_196);
  nand2 I005_214(w_005_214, w_003_050, w_004_319);
  nand2 I005_215(w_005_215, w_004_167, w_000_244);
  or2  I005_216(w_005_216, w_000_245, w_003_091);
  nand2 I005_217(w_005_217, w_003_012, w_001_004);
  or2  I005_218(w_005_218, w_003_096, w_003_041);
  not1 I005_219(w_005_219, w_003_021);
  and2 I005_220(w_005_220, w_003_023, w_001_001);
  nand2 I005_221(w_005_221, w_002_011, w_000_077);
  not1 I005_222(w_005_222, w_000_190);
  nand2 I005_223(w_005_223, w_003_030, w_002_002);
  nand2 I005_224(w_005_224, w_001_006, w_003_007);
  and2 I005_225(w_005_225, w_003_001, w_001_006);
  nand2 I005_226(w_005_226, w_004_418, w_001_006);
  nand2 I005_227(w_005_227, w_003_034, w_000_197);
  or2  I005_228(w_005_228, w_003_070, w_001_000);
  or2  I005_229(w_005_229, w_000_246, w_004_253);
  nand2 I005_230(w_005_230, w_001_006, w_004_301);
  nand2 I005_231(w_005_231, w_000_247, w_001_000);
  not1 I005_232(w_005_232, w_001_000);
  and2 I005_233(w_005_233, w_002_019, w_003_073);
  or2  I005_235(w_005_235, w_002_026, w_003_042);
  not1 I005_236(w_005_236, w_002_007);
  or2  I005_237(w_005_237, w_003_003, w_002_001);
  not1 I005_238(w_005_238, w_004_226);
  not1 I005_239(w_005_239, w_001_002);
  nand2 I005_241(w_005_241, w_002_001, w_004_464);
  and2 I005_242(w_005_242, w_000_066, w_000_250);
  and2 I005_243(w_005_243, w_004_020, w_002_005);
  or2  I005_244(w_005_244, w_002_008, w_000_251);
  nand2 I005_245(w_005_245, w_000_082, w_000_252);
  not1 I005_246(w_005_246, w_003_008);
  or2  I005_250(w_005_250, w_001_006, w_002_019);
  not1 I005_251(w_005_251, w_000_253);
  or2  I005_252(w_005_252, w_000_070, w_001_002);
  not1 I006_000(w_006_000, w_001_002);
  not1 I007_001(w_007_001, w_003_087);
  or2  I007_002(w_007_002, w_005_044, w_001_001);
  nand2 I007_003(w_007_003, w_004_280, w_000_254);
  not1 I007_004(w_007_004, w_000_255);
  and2 I007_005(w_007_005, w_000_181, w_005_050);
  or2  I007_006(w_007_006, w_006_000, w_001_004);
  and2 I007_007(w_007_007, w_006_000, w_002_011);
  not1 I007_008(w_007_008, w_003_037);
  nand2 I007_009(w_007_009, w_006_000, w_005_040);
  or2  I007_013(w_007_013, w_000_014, w_002_019);
  or2  I007_014(w_007_014, w_004_175, w_001_005);
  not1 I007_015(w_007_015, w_004_005);
  not1 I007_016(w_007_016, w_002_013);
  not1 I007_017(w_007_017, w_001_004);
  nand2 I007_018(w_007_018, w_005_015, w_004_172);
  nand2 I007_019(w_007_019, w_004_417, w_003_037);
  nand2 I007_020(w_007_020, w_001_002, w_004_124);
  nand2 I007_021(w_007_021, w_004_133, w_004_308);
  or2  I007_022(w_007_022, w_000_256, w_002_013);
  and2 I007_023(w_007_023, w_002_027, w_006_000);
  or2  I007_025(w_007_025, w_005_153, w_006_000);
  not1 I007_026(w_007_026, w_000_257);
  or2  I007_027(w_007_027, w_001_004, w_006_000);
  not1 I007_029(w_007_029, w_001_005);
  not1 I007_030(w_007_030, w_004_086);
  not1 I007_031(w_007_031, w_003_001);
  not1 I007_032(w_007_032, w_005_165);
  nand2 I007_033(w_007_033, w_003_076, w_000_189);
  and2 I007_035(w_007_035, w_001_005, w_000_258);
  not1 I007_038(w_007_038, w_006_000);
  or2  I007_039(w_007_039, w_003_078, w_000_235);
  or2  I007_040(w_007_040, w_004_072, w_004_192);
  not1 I007_041(w_007_041, w_002_004);
  not1 I007_042(w_007_042, w_002_027);
  nand2 I007_043(w_007_043, w_005_062, w_001_002);
  and2 I007_044(w_007_044, w_005_094, w_001_005);
  or2  I007_045(w_007_045, w_005_221, w_006_000);
  nand2 I007_046(w_007_046, w_002_003, w_001_004);
  and2 I007_047(w_007_047, w_003_099, w_004_388);
  nand2 I007_048(w_007_048, w_006_000, w_004_059);
  and2 I007_049(w_007_049, w_006_000, w_005_177);
  and2 I007_050(w_007_050, w_006_000, w_004_085);
  or2  I007_051(w_007_051, w_001_000, w_005_108);
  or2  I007_052(w_007_052, w_006_000, w_005_210);
  nand2 I007_053(w_007_053, w_006_000, w_002_014);
  or2  I007_055(w_007_055, w_002_017, w_003_023);
  or2  I007_056(w_007_056, w_004_384, w_002_003);
  or2  I007_057(w_007_057, w_006_000, w_000_190);
  or2  I007_058(w_007_058, w_003_051, w_005_155);
  not1 I007_059(w_007_059, w_000_206);
  and2 I007_060(w_007_060, w_002_001, w_003_048);
  nand2 I007_061(w_007_061, w_004_211, w_003_096);
  or2  I007_062(w_007_062, w_006_000, w_004_204);
  not1 I007_063(w_007_063, w_006_000);
  nand2 I007_064(w_007_064, w_003_040, w_001_002);
  or2  I007_065(w_007_065, w_002_004, w_001_001);
  not1 I007_066(w_007_066, w_002_010);
  not1 I007_068(w_007_068, w_002_011);
  and2 I007_069(w_007_069, w_000_260, w_005_193);
  or2  I007_070(w_007_070, w_004_324, w_003_096);
  nand2 I007_071(w_007_071, w_003_023, w_006_000);
  and2 I007_072(w_007_072, w_001_000, w_002_027);
  nand2 I007_073(w_007_073, w_004_094, w_000_102);
  and2 I007_074(w_007_074, w_001_000, w_002_027);
  and2 I007_075(w_007_075, w_003_050, w_002_027);
  not1 I007_076(w_007_076, w_004_114);
  not1 I007_077(w_007_077, w_000_261);
  not1 I007_078(w_007_078, w_003_096);
  or2  I007_080(w_007_080, w_005_037, w_005_184);
  and2 I007_081(w_007_081, w_001_000, w_001_002);
  and2 I007_082(w_007_082, w_002_013, w_001_004);
  or2  I007_083(w_007_083, w_005_200, w_006_000);
  nand2 I007_084(w_007_084, w_006_000, w_001_002);
  or2  I007_085(w_007_085, w_001_001, w_004_320);
  not1 I007_086(w_007_086, w_004_058);
  nand2 I007_087(w_007_087, w_000_095, w_000_262);
  and2 I007_088(w_007_088, w_006_000, w_004_427);
  not1 I007_089(w_007_089, w_003_065);
  nand2 I007_090(w_007_090, w_001_004, w_003_034);
  and2 I007_091(w_007_091, w_000_093, w_001_004);
  not1 I007_092(w_007_092, w_000_263);
  or2  I007_094(w_007_094, w_005_119, w_005_046);
  and2 I007_095(w_007_095, w_003_010, w_003_059);
  not1 I007_097(w_007_097, w_005_215);
  or2  I007_098(w_007_098, w_000_264, w_006_000);
  or2  I007_099(w_007_099, w_004_221, w_003_082);
  not1 I007_100(w_007_100, w_001_005);
  and2 I007_101(w_007_101, w_005_089, w_006_000);
  nand2 I007_104(w_007_104, w_006_000, w_000_265);
  not1 I007_105(w_007_105, w_000_149);
  nand2 I007_106(w_007_106, w_004_222, w_001_003);
  or2  I007_107(w_007_107, w_003_021, w_001_003);
  not1 I007_108(w_007_108, w_000_266);
  and2 I007_109(w_007_109, w_001_000, w_006_000);
  not1 I007_113(w_007_113, w_002_002);
  and2 I007_115(w_007_115, w_002_019, w_004_282);
  nand2 I007_116(w_007_116, w_006_000, w_003_082);
  not1 I007_117(w_007_117, w_005_207);
  or2  I007_118(w_007_118, w_003_086, w_005_005);
  or2  I007_119(w_007_119, w_004_104, w_005_236);
  not1 I007_120(w_007_120, w_005_067);
  and2 I007_121(w_007_121, w_006_000, w_003_042);
  and2 I007_122(w_007_122, w_003_046, w_005_058);
  or2  I007_123(w_007_123, w_002_025, w_001_000);
  nand2 I007_124(w_007_124, w_004_263, w_004_009);
  or2  I007_125(w_007_125, w_003_017, w_004_456);
  nand2 I007_126(w_007_126, w_002_018, w_002_016);
  or2  I007_128(w_007_128, w_004_228, w_004_318);
  not1 I007_129(w_007_129, w_003_024);
  or2  I007_131(w_007_131, w_005_156, w_002_005);
  or2  I007_134(w_007_134, w_004_349, w_005_225);
  not1 I007_135(w_007_135, w_001_002);
  and2 I007_136(w_007_136, w_002_017, w_001_003);
  or2  I007_137(w_007_137, w_004_029, w_000_093);
  not1 I007_138(w_007_138, w_005_101);
  nand2 I007_141(w_007_141, w_003_041, w_004_051);
  nand2 I007_142(w_007_142, w_005_109, w_001_002);
  not1 I007_143(w_007_143, w_002_014);
  nand2 I007_144(w_007_144, w_000_259, w_006_000);
  and2 I007_146(w_007_146, w_006_000, w_000_269);
  or2  I007_147(w_007_147, w_006_000, w_000_270);
  nand2 I007_148(w_007_148, w_004_467, w_002_020);
  and2 I007_154(w_007_154, w_006_000, w_004_357);
  and2 I007_156(w_007_156, w_003_091, w_004_321);
  or2  I007_159(w_007_159, w_005_216, w_006_000);
  or2  I007_160(w_007_160, w_003_079, w_005_227);
  nand2 I007_163(w_007_163, w_004_287, w_002_003);
  and2 I007_164(w_007_164, w_002_008, w_006_000);
  and2 I007_165(w_007_165, w_004_087, w_005_096);
  nand2 I007_166(w_007_166, w_004_325, w_002_011);
  and2 I007_167(w_007_167, w_000_272, w_002_013);
  nand2 I007_168(w_007_168, w_006_000, w_001_004);
  or2  I007_170(w_007_170, w_006_000, w_003_052);
  or2  I007_171(w_007_171, w_002_022, w_003_023);
  nand2 I007_172(w_007_172, w_000_273, w_000_008);
  or2  I007_173(w_007_173, w_002_003, w_003_000);
  and2 I007_174(w_007_174, w_000_110, w_004_429);
  not1 I007_175(w_007_175, w_004_297);
  and2 I007_176(w_007_176, w_001_004, w_002_026);
  not1 I007_177(w_007_177, w_005_033);
  nand2 I007_178(w_007_178, w_005_103, w_004_104);
  nand2 I007_180(w_007_180, w_000_274, w_006_000);
  nand2 I007_181(w_007_181, w_006_000, w_002_017);
  nand2 I007_182(w_007_182, w_004_222, w_001_006);
  nand2 I007_183(w_007_183, w_001_000, w_002_026);
  or2  I007_184(w_007_184, w_003_053, w_002_003);
  nand2 I007_186(w_007_186, w_005_004, w_001_004);
  nand2 I007_187(w_007_187, w_006_000, w_000_230);
  nand2 I007_188(w_007_188, w_006_000, w_001_004);
  or2  I007_189(w_007_189, w_002_001, w_006_000);
  and2 I007_190(w_007_190, w_004_005, w_005_122);
  nand2 I007_192(w_007_192, w_005_083, w_001_000);
  and2 I007_193(w_007_193, w_004_282, w_005_194);
  and2 I007_194(w_007_194, w_002_025, w_001_004);
  not1 I007_195(w_007_195, w_004_051);
  and2 I007_196(w_007_196, w_001_000, w_004_062);
  not1 I007_197(w_007_197, w_000_036);
  not1 I007_199(w_007_199, w_000_215);
  not1 I007_200(w_007_200, w_004_372);
  or2  I007_203(w_007_203, w_000_277, w_006_000);
  nand2 I007_204(w_007_204, w_001_006, w_005_187);
  nand2 I007_206(w_007_206, w_005_034, w_001_005);
  nand2 I007_208(w_007_208, w_000_061, w_005_216);
  not1 I007_209(w_007_209, w_005_024);
  nand2 I007_210(w_007_210, w_006_000, w_002_020);
  nand2 I007_211(w_007_211, w_002_013, w_000_279);
  or2  I007_213(w_007_213, w_001_003, w_002_003);
  not1 I007_214(w_007_214, w_003_073);
  nand2 I007_215(w_007_215, w_001_005, w_003_010);
  or2  I007_216(w_007_216, w_005_200, w_002_002);
  and2 I007_219(w_007_219, w_004_329, w_000_063);
  or2  I007_221(w_007_221, w_001_004, w_002_022);
  or2  I007_222(w_007_222, w_002_003, w_006_000);
  not1 I007_224(w_007_224, w_004_447);
  and2 I007_225(w_007_225, w_006_000, w_001_000);
  or2  I007_226(w_007_226, w_000_280, w_002_002);
  or2  I007_227(w_007_227, w_005_012, w_005_074);
  and2 I007_228(w_007_228, w_000_202, w_006_000);
  or2  I007_229(w_007_229, w_004_386, w_002_020);
  or2  I007_230(w_007_230, w_004_385, w_000_281);
  or2  I007_231(w_007_231, w_004_002, w_003_060);
  or2  I007_233(w_007_233, w_002_022, w_005_101);
  or2  I007_234(w_007_234, w_000_282, w_003_063);
  and2 I007_238(w_007_238, w_002_025, w_004_127);
  and2 I007_239(w_007_239, w_003_077, w_006_000);
  nand2 I007_240(w_007_240, w_001_001, w_004_031);
  nand2 I007_241(w_007_241, w_004_104, w_003_004);
  nand2 I007_242(w_007_242, w_000_035, w_004_441);
  nand2 I007_243(w_007_243, w_005_017, w_000_283);
  or2  I007_244(w_007_244, w_001_006, w_001_004);
  or2  I007_245(w_007_245, w_001_004, w_000_229);
  not1 I007_246(w_007_246, w_000_284);
  or2  I007_247(w_007_247, w_004_388, w_001_002);
  and2 I007_248(w_007_248, w_005_018, w_002_010);
  or2  I007_249(w_007_249, w_000_119, w_004_240);
  not1 I007_250(w_007_250, w_005_123);
  nand2 I007_251(w_007_251, w_004_431, w_000_102);
  and2 I007_252(w_007_252, w_006_000, w_004_088);
  or2  I007_253(w_007_253, w_004_445, w_000_285);
  not1 I007_254(w_007_254, w_000_155);
  not1 I007_255(w_007_255, w_003_071);
  not1 I007_258(w_007_258, w_006_000);
  not1 I007_259(w_007_259, w_005_231);
  or2  I007_260(w_007_260, w_005_086, w_001_000);
  or2  I007_261(w_007_261, w_005_173, w_005_158);
  not1 I007_262(w_007_262, w_006_000);
  and2 I007_263(w_007_263, w_006_000, w_004_201);
  or2  I007_264(w_007_264, w_000_144, w_005_151);
  nand2 I007_265(w_007_265, w_001_006, w_004_018);
  nand2 I007_266(w_007_266, w_000_002, w_002_005);
  or2  I007_267(w_007_267, w_003_036, w_005_003);
  nand2 I007_268(w_007_268, w_004_167, w_002_018);
  and2 I007_269(w_007_269, w_004_418, w_003_079);
  nand2 I007_270(w_007_270, w_005_190, w_004_070);
  or2  I007_271(w_007_271, w_003_006, w_005_243);
  and2 I007_272(w_007_272, w_005_023, w_003_002);
  or2  I007_273(w_007_273, w_006_000, w_004_094);
  not1 I007_275(w_007_275, w_005_036);
  nand2 I007_276(w_007_276, w_003_083, w_002_010);
  and2 I007_278(w_007_278, w_006_000, w_002_014);
  and2 I007_281(w_007_281, w_000_286, w_005_245);
  not1 I007_283(w_007_283, w_005_035);
  nand2 I007_284(w_007_284, w_002_024, w_006_000);
  or2  I007_285(w_007_285, w_002_021, w_005_154);
  nand2 I007_286(w_007_286, w_003_009, w_004_122);
  not1 I007_288(w_007_288, w_005_104);
  or2  I007_290(w_007_290, w_001_002, w_006_000);
  not1 I007_292(w_007_292, w_002_003);
  nand2 I007_293(w_007_293, w_005_227, w_002_010);
  and2 I007_296(w_007_296, w_004_164, w_006_000);
  nand2 I007_297(w_007_297, w_003_018, w_001_002);
  nand2 I007_298(w_007_298, w_001_002, w_003_060);
  and2 I007_299(w_007_299, w_002_021, w_006_000);
  and2 I007_300(w_007_300, w_006_000, w_002_023);
  nand2 I007_302(w_007_302, w_003_052, w_004_253);
  not1 I007_303(w_007_303, w_005_027);
  nand2 I007_305(w_007_305, w_001_004, w_004_289);
  and2 I007_306(w_007_306, w_002_012, w_001_001);
  and2 I007_307(w_007_307, w_003_079, w_003_076);
  and2 I007_308(w_007_308, w_001_005, w_005_147);
  and2 I007_309(w_007_309, w_003_048, w_001_000);
  or2  I007_314(w_007_314, w_001_001, w_001_003);
  nand2 I007_315(w_007_315, w_006_000, w_003_029);
  nand2 I007_316(w_007_316, w_004_204, w_006_000);
  not1 I007_317(w_007_317, w_003_054);
  nand2 I007_319(w_007_319, w_000_291, w_004_401);
  or2  I007_320(w_007_320, w_003_030, w_005_022);
  not1 I007_321(w_007_321, w_004_024);
  or2  I007_322(w_007_322, w_001_005, w_000_104);
  nand2 I007_324(w_007_324, w_003_093, w_005_216);
  nand2 I007_325(w_007_325, w_002_022, w_000_163);
  or2  I007_328(w_007_328, w_001_003, w_000_292);
  not1 I007_329(w_007_329, w_002_012);
  not1 I007_333(w_007_333, w_006_000);
  or2  I007_337(w_007_337, w_004_060, w_000_294);
  nand2 I007_340(w_007_340, w_006_000, w_004_358);
  and2 I007_341(w_007_341, w_006_000, w_000_295);
  and2 I007_342(w_007_342, w_003_075, w_001_004);
  and2 I007_343(w_007_343, w_003_037, w_002_014);
  and2 I007_344(w_007_344, w_004_234, w_000_296);
  nand2 I007_345(w_007_345, w_004_234, w_000_297);
  and2 I007_347(w_007_347, w_002_013, w_006_000);
  and2 I007_348(w_007_348, w_006_000, w_004_340);
  not1 I007_349(w_007_349, w_004_131);
  nand2 I007_350(w_007_350, w_000_298, w_004_224);
  not1 I007_352(w_007_352, w_003_032);
  and2 I007_354(w_007_354, w_001_001, w_003_096);
  not1 I007_355(w_007_355, w_001_003);
  not1 I007_356(w_007_356, w_002_023);
  not1 I007_357(w_007_357, w_001_001);
  or2  I007_359(w_007_359, w_000_300, w_005_196);
  not1 I007_360(w_007_360, w_000_113);
  and2 I007_361(w_007_361, w_000_270, w_003_056);
  nand2 I007_362(w_007_362, w_003_054, w_004_127);
  and2 I007_363(w_007_363, w_002_025, w_005_104);
  nand2 I007_364(w_007_364, w_006_000, w_005_093);
  nand2 I007_366(w_007_366, w_006_000, w_002_008);
  or2  I007_367(w_007_367, w_006_000, w_002_021);
  and2 I007_368(w_007_368, w_001_006, w_001_000);
  not1 I007_370(w_007_370, w_003_099);
  or2  I007_371(w_007_371, w_002_004, w_001_000);
  or2  I007_372(w_007_372, w_001_002, w_005_088);
  and2 I007_373(w_007_373, w_000_181, w_001_000);
  or2  I007_374(w_007_374, w_001_000, w_005_142);
  and2 I007_376(w_007_376, w_006_000, w_002_000);
  and2 I007_377(w_007_377, w_001_004, w_005_037);
  nand2 I007_378(w_007_378, w_001_002, w_004_327);
  nand2 I007_379(w_007_379, w_000_072, w_004_234);
  or2  I007_380(w_007_380, w_006_000, w_003_092);
  and2 I007_381(w_007_381, w_004_152, w_002_004);
  nand2 I007_382(w_007_382, w_005_095, w_005_231);
  nand2 I007_383(w_007_383, w_000_302, w_006_000);
  and2 I007_385(w_007_385, w_005_065, w_006_000);
  nand2 I007_386(w_007_386, w_003_071, w_000_167);
  not1 I007_388(w_007_388, w_000_303);
  nand2 I007_389(w_007_389, w_003_068, w_005_162);
  nand2 I007_390(w_007_390, w_001_005, w_001_004);
  nand2 I007_391(w_007_391, w_004_319, w_005_113);
  or2  I007_394(w_007_394, w_004_080, w_004_303);
  not1 I007_396(w_007_396, w_000_039);
  or2  I007_398(w_007_398, w_000_305, w_002_013);
  and2 I007_400(w_007_400, w_006_000, w_000_306);
  or2  I007_403(w_007_403, w_005_095, w_006_000);
  not1 I007_404(w_007_404, w_005_082);
  not1 I008_000(w_008_000, w_001_004);
  nand2 I008_001(w_008_001, w_000_307, w_000_073);
  nand2 I008_003(w_008_003, w_002_001, w_007_077);
  nand2 I008_004(w_008_004, w_007_039, w_005_094);
  not1 I008_005(w_008_005, w_006_000);
  or2  I008_008(w_008_008, w_007_377, w_005_163);
  not1 I008_010(w_008_010, w_001_000);
  or2  I008_011(w_008_011, w_000_203, w_006_000);
  or2  I008_012(w_008_012, w_004_032, w_007_124);
  or2  I008_013(w_008_013, w_004_143, w_005_141);
  or2  I008_014(w_008_014, w_002_005, w_006_000);
  or2  I008_015(w_008_015, w_003_065, w_000_308);
  not1 I008_016(w_008_016, w_001_002);
  and2 I008_017(w_008_017, w_002_001, w_005_138);
  or2  I008_018(w_008_018, w_003_009, w_006_000);
  nand2 I008_020(w_008_020, w_004_184, w_000_234);
  not1 I008_022(w_008_022, w_003_033);
  and2 I008_023(w_008_023, w_004_398, w_004_223);
  nand2 I008_024(w_008_024, w_001_004, w_004_348);
  nand2 I008_025(w_008_025, w_003_007, w_004_189);
  nand2 I008_026(w_008_026, w_003_071, w_006_000);
  nand2 I008_027(w_008_027, w_006_000, w_004_432);
  not1 I008_028(w_008_028, w_007_084);
  and2 I008_029(w_008_029, w_002_013, w_004_427);
  nand2 I008_030(w_008_030, w_000_150, w_006_000);
  nand2 I008_031(w_008_031, w_003_039, w_006_000);
  or2  I008_032(w_008_032, w_003_073, w_000_162);
  not1 I008_033(w_008_033, w_006_000);
  or2  I008_034(w_008_034, w_004_351, w_005_112);
  not1 I008_035(w_008_035, w_005_200);
  nand2 I008_037(w_008_037, w_006_000, w_007_376);
  and2 I008_038(w_008_038, w_001_001, w_007_394);
  not1 I008_039(w_008_039, w_005_050);
  or2  I008_040(w_008_040, w_004_023, w_004_098);
  or2  I008_041(w_008_041, w_002_007, w_001_004);
  or2  I008_043(w_008_043, w_005_130, w_003_040);
  and2 I008_045(w_008_045, w_002_023, w_003_034);
  nand2 I008_046(w_008_046, w_003_098, w_005_207);
  not1 I008_047(w_008_047, w_004_234);
  nand2 I008_048(w_008_048, w_000_309, w_007_290);
  and2 I008_050(w_008_050, w_002_014, w_003_092);
  not1 I008_051(w_008_051, w_002_004);
  not1 I008_052(w_008_052, w_000_310);
  or2  I008_053(w_008_053, w_003_075, w_001_004);
  not1 I008_054(w_008_054, w_005_138);
  nand2 I008_056(w_008_056, w_004_353, w_005_074);
  not1 I008_057(w_008_057, w_000_311);
  and2 I008_058(w_008_058, w_003_056, w_003_037);
  and2 I008_059(w_008_059, w_007_240, w_004_347);
  or2  I008_060(w_008_060, w_007_017, w_002_017);
  or2  I008_061(w_008_061, w_007_160, w_000_302);
  nand2 I008_062(w_008_062, w_001_005, w_006_000);
  not1 I008_063(w_008_063, w_004_452);
  and2 I008_064(w_008_064, w_004_323, w_005_107);
  or2  I008_065(w_008_065, w_000_201, w_001_004);
  or2  I008_066(w_008_066, w_005_046, w_002_004);
  and2 I008_067(w_008_067, w_004_053, w_001_004);
  or2  I008_068(w_008_068, w_001_005, w_000_026);
  and2 I008_070(w_008_070, w_004_307, w_000_257);
  and2 I008_072(w_008_072, w_001_004, w_006_000);
  or2  I008_073(w_008_073, w_006_000, w_002_000);
  or2  I008_074(w_008_074, w_007_083, w_004_156);
  nand2 I008_075(w_008_075, w_004_136, w_006_000);
  and2 I008_076(w_008_076, w_006_000, w_005_165);
  not1 I008_077(w_008_077, w_006_000);
  or2  I008_078(w_008_078, w_006_000, w_001_006);
  or2  I008_079(w_008_079, w_002_010, w_000_193);
  not1 I008_080(w_008_080, w_002_025);
  and2 I008_081(w_008_081, w_001_005, w_000_313);
  or2  I008_082(w_008_082, w_004_465, w_003_092);
  or2  I008_083(w_008_083, w_001_004, w_006_000);
  nand2 I008_084(w_008_084, w_004_431, w_000_314);
  or2  I008_085(w_008_085, w_001_002, w_002_020);
  or2  I008_086(w_008_086, w_002_009, w_003_006);
  not1 I008_087(w_008_087, w_007_080);
  nand2 I008_088(w_008_088, w_007_315, w_000_039);
  and2 I008_089(w_008_089, w_004_336, w_002_021);
  or2  I008_090(w_008_090, w_000_108, w_000_093);
  nand2 I008_091(w_008_091, w_000_315, w_001_004);
  not1 I008_092(w_008_092, w_003_095);
  nand2 I008_093(w_008_093, w_006_000, w_002_022);
  nand2 I008_095(w_008_095, w_000_273, w_003_022);
  or2  I008_096(w_008_096, w_005_033, w_002_018);
  or2  I008_098(w_008_098, w_002_002, w_006_000);
  and2 I008_099(w_008_099, w_002_009, w_007_160);
  nand2 I008_100(w_008_100, w_002_006, w_000_236);
  or2  I008_102(w_008_102, w_000_242, w_001_001);
  nand2 I008_103(w_008_103, w_006_000, w_001_001);
  or2  I008_104(w_008_104, w_003_001, w_002_017);
  not1 I008_105(w_008_105, w_001_006);
  not1 I008_106(w_008_106, w_003_064);
  not1 I008_107(w_008_107, w_003_079);
  or2  I008_109(w_008_109, w_005_196, w_006_000);
  not1 I008_110(w_008_110, w_003_013);
  or2  I008_111(w_008_111, w_002_001, w_001_000);
  and2 I008_112(w_008_112, w_001_002, w_002_023);
  not1 I008_113(w_008_113, w_003_063);
  or2  I008_114(w_008_114, w_005_134, w_000_317);
  nand2 I008_115(w_008_115, w_006_000, w_003_044);
  or2  I008_116(w_008_116, w_001_004, w_003_031);
  not1 I008_117(w_008_117, w_006_000);
  nand2 I008_118(w_008_118, w_000_105, w_000_003);
  not1 I008_119(w_008_119, w_001_005);
  and2 I008_120(w_008_120, w_004_027, w_003_098);
  or2  I008_121(w_008_121, w_000_318, w_001_001);
  and2 I008_123(w_008_123, w_001_005, w_003_002);
  nand2 I008_124(w_008_124, w_002_019, w_002_014);
  and2 I008_125(w_008_125, w_002_010, w_002_024);
  nand2 I008_126(w_008_126, w_002_004, w_006_000);
  not1 I008_127(w_008_127, w_007_325);
  and2 I008_128(w_008_128, w_001_001, w_001_006);
  not1 I008_130(w_008_130, w_003_053);
  not1 I008_131(w_008_131, w_005_038);
  and2 I008_132(w_008_132, w_000_319, w_002_017);
  not1 I008_133(w_008_133, w_004_015);
  not1 I008_134(w_008_134, w_007_098);
  nand2 I008_135(w_008_135, w_006_000, w_005_008);
  nand2 I008_137(w_008_137, w_007_007, w_005_154);
  nand2 I008_138(w_008_138, w_004_100, w_004_342);
  and2 I008_139(w_008_139, w_005_090, w_002_014);
  and2 I008_140(w_008_140, w_007_085, w_003_042);
  not1 I008_142(w_008_142, w_000_205);
  and2 I008_143(w_008_143, w_005_114, w_007_071);
  not1 I008_145(w_008_145, w_007_322);
  not1 I008_146(w_008_146, w_004_412);
  and2 I008_148(w_008_148, w_006_000, w_002_027);
  not1 I008_149(w_008_149, w_005_184);
  not1 I008_150(w_008_150, w_002_025);
  or2  I008_152(w_008_152, w_006_000, w_002_004);
  nand2 I008_153(w_008_153, w_000_219, w_003_049);
  and2 I008_154(w_008_154, w_001_005, w_004_009);
  and2 I008_156(w_008_156, w_005_157, w_005_009);
  nand2 I008_157(w_008_157, w_000_320, w_002_002);
  and2 I008_161(w_008_161, w_007_259, w_002_002);
  not1 I008_162(w_008_162, w_002_023);
  nand2 I008_165(w_008_165, w_004_413, w_005_104);
  and2 I008_166(w_008_166, w_006_000, w_007_131);
  or2  I008_168(w_008_168, w_003_046, w_007_181);
  and2 I008_169(w_008_169, w_001_000, w_004_000);
  nand2 I008_173(w_008_173, w_003_098, w_002_018);
  not1 I008_175(w_008_175, w_005_236);
  or2  I008_176(w_008_176, w_003_003, w_002_020);
  and2 I008_177(w_008_177, w_006_000, w_000_321);
  or2  I008_179(w_008_179, w_000_322, w_002_026);
  nand2 I008_180(w_008_180, w_005_244, w_001_005);
  or2  I008_183(w_008_183, w_004_317, w_001_004);
  or2  I008_184(w_008_184, w_001_003, w_002_014);
  or2  I008_185(w_008_185, w_000_323, w_002_021);
  and2 I008_186(w_008_186, w_004_020, w_000_133);
  and2 I008_187(w_008_187, w_001_002, w_000_324);
  or2  I008_190(w_008_190, w_006_000, w_002_004);
  nand2 I008_191(w_008_191, w_004_011, w_005_169);
  not1 I008_193(w_008_193, w_004_465);
  and2 I008_195(w_008_195, w_006_000, w_005_127);
  nand2 I008_196(w_008_196, w_004_181, w_007_188);
  or2  I008_198(w_008_198, w_003_084, w_001_003);
  and2 I008_199(w_008_199, w_003_048, w_005_184);
  nand2 I008_200(w_008_200, w_003_015, w_003_049);
  not1 I008_201(w_008_201, w_001_001);
  not1 I008_202(w_008_202, w_007_241);
  nand2 I008_203(w_008_203, w_007_192, w_000_325);
  and2 I008_205(w_008_205, w_003_100, w_001_002);
  not1 I008_206(w_008_206, w_004_154);
  and2 I008_207(w_008_207, w_005_062, w_007_272);
  or2  I008_208(w_008_208, w_000_328, w_002_019);
  and2 I008_209(w_008_209, w_001_004, w_004_293);
  or2  I008_210(w_008_210, w_004_265, w_001_002);
  and2 I008_212(w_008_212, w_005_050, w_003_043);
  not1 I008_215(w_008_215, w_006_000);
  nand2 I008_216(w_008_216, w_002_018, w_000_134);
  or2  I008_218(w_008_218, w_004_374, w_005_106);
  or2  I008_219(w_008_219, w_000_103, w_003_033);
  not1 I008_223(w_008_223, w_002_016);
  and2 I008_225(w_008_225, w_002_020, w_001_005);
  or2  I008_226(w_008_226, w_002_003, w_000_129);
  and2 I008_228(w_008_228, w_001_000, w_004_333);
  and2 I008_230(w_008_230, w_001_000, w_007_394);
  not1 I008_231(w_008_231, w_003_032);
  nand2 I008_233(w_008_233, w_007_180, w_004_004);
  or2  I008_234(w_008_234, w_007_076, w_004_417);
  and2 I008_236(w_008_236, w_007_190, w_000_200);
  nand2 I008_237(w_008_237, w_001_004, w_006_000);
  not1 I008_238(w_008_238, w_002_016);
  and2 I008_239(w_008_239, w_007_136, w_000_090);
  and2 I008_240(w_008_240, w_004_094, w_006_000);
  not1 I008_241(w_008_241, w_002_004);
  nand2 I008_242(w_008_242, w_007_195, w_003_095);
  and2 I008_243(w_008_243, w_002_024, w_000_130);
  nand2 I008_244(w_008_244, w_001_001, w_005_039);
  or2  I008_245(w_008_245, w_007_300, w_002_006);
  or2  I008_246(w_008_246, w_002_004, w_005_045);
  not1 I008_250(w_008_250, w_005_085);
  or2  I008_251(w_008_251, w_006_000, w_001_002);
  nand2 I008_252(w_008_252, w_003_014, w_004_257);
  or2  I008_253(w_008_253, w_001_006, w_004_277);
  and2 I008_254(w_008_254, w_005_190, w_006_000);
  nand2 I008_255(w_008_255, w_003_030, w_001_000);
  and2 I008_256(w_008_256, w_003_037, w_001_005);
  and2 I008_258(w_008_258, w_000_331, w_005_087);
  nand2 I008_260(w_008_260, w_000_332, w_005_117);
  or2  I008_261(w_008_261, w_004_057, w_003_095);
  and2 I008_263(w_008_263, w_001_006, w_007_021);
  not1 I008_264(w_008_264, w_007_015);
  nand2 I008_268(w_008_268, w_001_002, w_004_065);
  and2 I008_269(w_008_269, w_002_022, w_005_219);
  or2  I008_270(w_008_270, w_004_022, w_007_251);
  and2 I008_271(w_008_271, w_000_335, w_000_336);
  nand2 I008_273(w_008_273, w_006_000, w_003_046);
  not1 I008_274(w_008_274, w_000_246);
  or2  I008_275(w_008_275, w_001_000, w_001_002);
  nand2 I008_276(w_008_276, w_003_083, w_004_410);
  not1 I008_277(w_008_277, w_000_260);
  not1 I008_280(w_008_280, w_006_000);
  and2 I008_282(w_008_282, w_006_000, w_002_007);
  not1 I008_283(w_008_283, w_001_000);
  not1 I008_287(w_008_287, w_001_005);
  or2  I008_288(w_008_288, w_006_000, w_001_002);
  and2 I008_290(w_008_290, w_002_008, w_005_194);
  or2  I008_291(w_008_291, w_005_019, w_006_000);
  nand2 I008_292(w_008_292, w_006_000, w_002_024);
  nand2 I008_294(w_008_294, w_001_005, w_000_338);
  nand2 I008_296(w_008_296, w_000_155, w_004_225);
  not1 I008_297(w_008_297, w_001_005);
  or2  I008_299(w_008_299, w_006_000, w_003_074);
  nand2 I008_300(w_008_300, w_005_107, w_007_314);
  not1 I008_302(w_008_302, w_007_051);
  nand2 I008_304(w_008_304, w_003_033, w_000_038);
  or2  I008_307(w_008_307, w_004_237, w_002_023);
  and2 I008_309(w_008_309, w_007_350, w_004_435);
  or2  I008_310(w_008_310, w_004_278, w_000_332);
  not1 I008_311(w_008_311, w_001_005);
  not1 I008_312(w_008_312, w_004_338);
  and2 I008_315(w_008_315, w_004_111, w_005_070);
  not1 I008_317(w_008_317, w_001_004);
  not1 I008_318(w_008_318, w_004_053);
  and2 I008_320(w_008_320, w_004_086, w_003_027);
  nand2 I008_321(w_008_321, w_003_061, w_001_000);
  not1 I008_324(w_008_324, w_003_075);
  and2 I008_325(w_008_325, w_003_037, w_004_001);
  or2  I008_327(w_008_327, w_003_021, w_000_027);
  not1 I008_329(w_008_329, w_006_000);
  not1 I008_331(w_008_331, w_002_021);
  or2  I008_333(w_008_333, w_005_034, w_003_043);
  and2 I008_337(w_008_337, w_007_199, w_002_022);
  and2 I008_342(w_008_342, w_006_000, w_002_018);
  and2 I008_343(w_008_343, w_007_070, w_003_059);
  nand2 I008_345(w_008_345, w_006_000, w_000_285);
  and2 I009_000(w_009_000, w_007_211, w_005_040);
  not1 I009_001(w_009_001, w_006_000);
  not1 I009_002(w_009_002, w_008_304);
  and2 I009_003(w_009_003, w_008_145, w_004_206);
  not1 I009_004(w_009_004, w_000_069);
  nand2 I009_005(w_009_005, w_005_133, w_005_046);
  nand2 I009_006(w_009_006, w_007_224, w_002_000);
  or2  I009_007(w_009_007, w_006_000, w_000_342);
  or2  I009_008(w_009_008, w_002_013, w_000_192);
  nand2 I009_009(w_009_009, w_006_000, w_008_288);
  and2 I009_010(w_009_010, w_001_004, w_001_000);
  nand2 I009_011(w_009_011, w_002_021, w_005_093);
  nand2 I009_012(w_009_012, w_002_009, w_008_073);
  not1 I009_013(w_009_013, w_001_005);
  nand2 I009_014(w_009_014, w_002_009, w_005_081);
  not1 I009_015(w_009_015, w_005_126);
  or2  I009_016(w_009_016, w_001_006, w_004_210);
  nand2 I009_017(w_009_017, w_005_057, w_005_179);
  and2 I009_018(w_009_018, w_007_226, w_004_007);
  or2  I009_019(w_009_019, w_006_000, w_003_073);
  nand2 I009_020(w_009_020, w_002_006, w_006_000);
  nand2 I009_021(w_009_021, w_002_024, w_008_145);
  not1 I009_022(w_009_022, w_004_067);
  nand2 I009_024(w_009_024, w_004_381, w_007_159);
  nand2 I009_025(w_009_025, w_000_166, w_007_345);
  nand2 I009_026(w_009_026, w_001_000, w_003_069);
  not1 I009_027(w_009_027, w_000_343);
  or2  I009_028(w_009_028, w_000_049, w_005_072);
  nand2 I009_029(w_009_029, w_008_145, w_005_096);
  or2  I009_030(w_009_030, w_004_297, w_008_059);
  not1 I009_031(w_009_031, w_007_064);
  or2  I009_032(w_009_032, w_007_231, w_005_197);
  not1 I009_033(w_009_033, w_004_274);
  or2  I009_034(w_009_034, w_006_000, w_002_000);
  not1 I009_035(w_009_035, w_003_041);
  and2 I009_036(w_009_036, w_005_225, w_007_107);
  or2  I009_037(w_009_037, w_002_005, w_005_220);
  or2  I009_038(w_009_038, w_002_018, w_001_002);
  or2  I009_040(w_009_040, w_006_000, w_003_086);
  not1 I009_041(w_009_041, w_004_384);
  and2 I009_042(w_009_042, w_007_129, w_000_344);
  not1 I009_043(w_009_043, w_006_000);
  and2 I009_044(w_009_044, w_008_236, w_004_148);
  not1 I009_045(w_009_045, w_004_251);
  nand2 I009_046(w_009_046, w_002_027, w_007_400);
  or2  I009_047(w_009_047, w_007_214, w_005_042);
  and2 I009_048(w_009_048, w_007_039, w_004_018);
  and2 I009_049(w_009_049, w_000_000, w_007_260);
  not1 I009_050(w_009_050, w_004_268);
  not1 I009_051(w_009_051, w_001_006);
  and2 I009_052(w_009_052, w_000_130, w_006_000);
  nand2 I009_054(w_009_054, w_008_343, w_006_000);
  nand2 I009_056(w_009_056, w_005_180, w_008_238);
  nand2 I009_058(w_009_058, w_004_260, w_005_031);
  nand2 I009_059(w_009_059, w_000_174, w_003_085);
  nand2 I009_061(w_009_061, w_006_000, w_005_013);
  nand2 I009_062(w_009_062, w_004_103, w_008_032);
  not1 I009_063(w_009_063, w_000_168);
  nand2 I009_064(w_009_064, w_003_072, w_000_016);
  or2  I009_065(w_009_065, w_003_047, w_005_136);
  not1 I009_067(w_009_067, w_001_006);
  nand2 I009_072(w_009_072, w_000_262, w_008_113);
  not1 I009_073(w_009_073, w_006_000);
  not1 I009_074(w_009_074, w_002_022);
  and2 I009_075(w_009_075, w_008_102, w_000_247);
  nand2 I009_076(w_009_076, w_005_085, w_000_346);
  and2 I009_077(w_009_077, w_007_319, w_008_051);
  nand2 I009_078(w_009_078, w_008_062, w_005_213);
  nand2 I009_079(w_009_079, w_006_000, w_000_176);
  not1 I009_080(w_009_080, w_007_008);
  and2 I009_081(w_009_081, w_007_030, w_006_000);
  or2  I009_083(w_009_083, w_005_023, w_002_009);
  not1 I009_084(w_009_084, w_008_116);
  or2  I009_086(w_009_086, w_006_000, w_003_031);
  and2 I009_088(w_009_088, w_004_239, w_007_367);
  nand2 I009_089(w_009_089, w_005_022, w_006_000);
  or2  I009_090(w_009_090, w_006_000, w_001_002);
  nand2 I009_091(w_009_091, w_008_093, w_001_005);
  or2  I009_092(w_009_092, w_003_072, w_004_311);
  or2  I009_093(w_009_093, w_006_000, w_004_112);
  or2  I009_094(w_009_094, w_008_104, w_003_083);
  and2 I009_096(w_009_096, w_005_218, w_005_039);
  and2 I009_098(w_009_098, w_001_006, w_007_154);
  or2  I009_099(w_009_099, w_005_163, w_006_000);
  not1 I009_101(w_009_101, w_006_000);
  not1 I009_103(w_009_103, w_000_347);
  nand2 I009_104(w_009_104, w_004_199, w_000_237);
  not1 I009_105(w_009_105, w_006_000);
  not1 I009_106(w_009_106, w_002_017);
  and2 I009_107(w_009_107, w_004_001, w_007_025);
  and2 I009_108(w_009_108, w_006_000, w_001_004);
  and2 I009_109(w_009_109, w_003_086, w_004_304);
  or2  I009_111(w_009_111, w_002_025, w_003_054);
  nand2 I009_112(w_009_112, w_007_108, w_006_000);
  or2  I009_113(w_009_113, w_004_188, w_008_008);
  and2 I009_115(w_009_115, w_004_245, w_008_090);
  nand2 I009_116(w_009_116, w_004_246, w_003_090);
  or2  I009_117(w_009_117, w_002_012, w_008_268);
  or2  I009_118(w_009_118, w_002_015, w_004_462);
  not1 I009_120(w_009_120, w_001_005);
  and2 I009_121(w_009_121, w_004_183, w_005_094);
  or2  I009_122(w_009_122, w_003_082, w_005_126);
  nand2 I009_123(w_009_123, w_008_025, w_004_291);
  or2  I009_124(w_009_124, w_003_059, w_006_000);
  not1 I009_125(w_009_125, w_001_002);
  not1 I009_126(w_009_126, w_001_001);
  nand2 I009_127(w_009_127, w_003_068, w_007_258);
  and2 I009_128(w_009_128, w_000_294, w_007_039);
  nand2 I009_129(w_009_129, w_008_135, w_007_352);
  and2 I009_130(w_009_130, w_007_229, w_008_022);
  not1 I009_131(w_009_131, w_002_025);
  or2  I009_132(w_009_132, w_004_316, w_002_009);
  not1 I009_133(w_009_133, w_001_002);
  or2  I009_134(w_009_134, w_002_007, w_000_348);
  nand2 I009_135(w_009_135, w_007_077, w_001_004);
  and2 I009_136(w_009_136, w_001_005, w_004_361);
  nand2 I009_137(w_009_137, w_000_091, w_006_000);
  not1 I009_139(w_009_139, w_007_343);
  and2 I009_140(w_009_140, w_006_000, w_001_000);
  not1 I009_142(w_009_142, w_002_001);
  not1 I009_143(w_009_143, w_001_006);
  or2  I009_144(w_009_144, w_004_372, w_006_000);
  and2 I009_145(w_009_145, w_002_023, w_004_190);
  or2  I009_146(w_009_146, w_006_000, w_005_096);
  and2 I009_147(w_009_147, w_001_004, w_007_144);
  and2 I009_148(w_009_148, w_006_000, w_002_008);
  nand2 I009_149(w_009_149, w_005_092, w_000_070);
  nand2 I009_151(w_009_151, w_001_003, w_001_006);
  nand2 I009_152(w_009_152, w_000_234, w_006_000);
  and2 I009_153(w_009_153, w_005_163, w_003_011);
  not1 I009_154(w_009_154, w_004_134);
  and2 I009_155(w_009_155, w_006_000, w_004_249);
  and2 I009_156(w_009_156, w_002_004, w_000_183);
  not1 I009_157(w_009_157, w_007_008);
  or2  I009_158(w_009_158, w_007_033, w_000_349);
  or2  I009_159(w_009_159, w_007_138, w_001_006);
  nand2 I009_160(w_009_160, w_005_098, w_008_239);
  not1 I009_161(w_009_161, w_004_373);
  not1 I009_162(w_009_162, w_008_090);
  or2  I009_163(w_009_163, w_007_196, w_004_463);
  and2 I009_164(w_009_164, w_003_053, w_004_307);
  nand2 I009_165(w_009_165, w_002_014, w_007_315);
  or2  I009_167(w_009_167, w_004_026, w_003_087);
  and2 I009_168(w_009_168, w_007_267, w_007_403);
  nand2 I009_169(w_009_169, w_000_194, w_008_001);
  or2  I009_170(w_009_170, w_005_245, w_007_216);
  not1 I009_171(w_009_171, w_005_227);
  and2 I009_172(w_009_172, w_001_000, w_006_000);
  or2  I009_173(w_009_173, w_007_357, w_007_361);
  nand2 I009_174(w_009_174, w_002_003, w_002_008);
  not1 I009_175(w_009_175, w_000_350);
  or2  I009_176(w_009_176, w_007_105, w_003_071);
  not1 I009_177(w_009_177, w_006_000);
  or2  I009_178(w_009_178, w_006_000, w_005_066);
  nand2 I009_179(w_009_179, w_005_214, w_002_016);
  and2 I009_181(w_009_181, w_001_003, w_008_206);
  nand2 I009_183(w_009_183, w_002_007, w_002_001);
  and2 I009_185(w_009_185, w_008_023, w_008_039);
  and2 I009_186(w_009_186, w_001_003, w_007_154);
  or2  I009_187(w_009_187, w_003_046, w_007_261);
  not1 I009_189(w_009_189, w_007_049);
  not1 I009_190(w_009_190, w_007_050);
  nand2 I009_191(w_009_191, w_000_351, w_001_001);
  nand2 I009_192(w_009_192, w_007_206, w_005_117);
  not1 I009_193(w_009_193, w_006_000);
  and2 I009_194(w_009_194, w_007_293, w_006_000);
  nand2 I009_196(w_009_196, w_002_012, w_007_344);
  or2  I009_197(w_009_197, w_001_003, w_004_187);
  or2  I009_198(w_009_198, w_003_022, w_004_252);
  or2  I009_199(w_009_199, w_003_004, w_005_094);
  or2  I009_200(w_009_200, w_000_282, w_000_340);
  and2 I009_202(w_009_202, w_003_082, w_007_023);
  and2 I009_203(w_009_203, w_002_009, w_008_001);
  and2 I009_204(w_009_204, w_004_070, w_008_175);
  or2  I009_206(w_009_206, w_002_018, w_007_081);
  and2 I009_208(w_009_208, w_002_020, w_004_472);
  and2 I009_209(w_009_209, w_002_000, w_004_031);
  nand2 I009_211(w_009_211, w_006_000, w_007_026);
  and2 I009_212(w_009_212, w_008_312, w_007_049);
  nand2 I009_213(w_009_213, w_007_100, w_008_107);
  nand2 I009_216(w_009_216, w_000_314, w_008_095);
  and2 I009_217(w_009_217, w_003_072, w_000_323);
  and2 I009_218(w_009_218, w_007_204, w_007_038);
  nand2 I009_220(w_009_220, w_003_080, w_002_010);
  and2 I009_221(w_009_221, w_006_000, w_005_021);
  not1 I009_222(w_009_222, w_007_032);
  and2 I009_223(w_009_223, w_007_385, w_005_158);
  or2  I009_224(w_009_224, w_006_000, w_002_015);
  nand2 I009_225(w_009_225, w_000_042, w_004_308);
  not1 I009_226(w_009_226, w_002_026);
  or2  I009_227(w_009_227, w_006_000, w_000_228);
  and2 I009_228(w_009_228, w_006_000, w_002_000);
  and2 I009_229(w_009_229, w_005_017, w_006_000);
  and2 I009_231(w_009_231, w_003_012, w_000_352);
  and2 I009_232(w_009_232, w_003_025, w_003_064);
  nand2 I009_233(w_009_233, w_007_056, w_006_000);
  not1 I009_234(w_009_234, w_004_227);
  or2  I009_235(w_009_235, w_004_451, w_006_000);
  or2  I009_236(w_009_236, w_003_063, w_008_234);
  and2 I009_237(w_009_237, w_007_379, w_006_000);
  or2  I010_002(w_010_002, w_004_325, w_004_241);
  or2  I010_004(w_010_004, w_008_033, w_001_004);
  or2  I010_005(w_010_005, w_003_086, w_005_125);
  and2 I010_007(w_010_007, w_005_245, w_002_009);
  and2 I010_008(w_010_008, w_001_002, w_009_075);
  and2 I010_009(w_010_009, w_002_013, w_008_105);
  not1 I010_012(w_010_012, w_006_000);
  or2  I010_013(w_010_013, w_002_013, w_007_267);
  not1 I010_014(w_010_014, w_009_206);
  not1 I010_015(w_010_015, w_002_023);
  nand2 I010_016(w_010_016, w_008_271, w_006_000);
  nand2 I010_018(w_010_018, w_005_019, w_001_003);
  nand2 I010_020(w_010_020, w_008_100, w_006_000);
  and2 I010_021(w_010_021, w_008_126, w_008_110);
  and2 I010_023(w_010_023, w_001_001, w_007_329);
  nand2 I010_024(w_010_024, w_008_050, w_007_199);
  nand2 I010_025(w_010_025, w_007_187, w_007_382);
  and2 I010_026(w_010_026, w_008_290, w_007_092);
  not1 I010_027(w_010_027, w_003_083);
  not1 I010_028(w_010_028, w_004_147);
  or2  I010_029(w_010_029, w_008_114, w_002_018);
  and2 I010_030(w_010_030, w_005_225, w_005_196);
  and2 I010_033(w_010_033, w_008_124, w_003_035);
  not1 I010_034(w_010_034, w_009_220);
  and2 I010_035(w_010_035, w_003_015, w_005_020);
  nand2 I010_036(w_010_036, w_008_183, w_007_033);
  and2 I010_037(w_010_037, w_004_230, w_001_006);
  not1 I010_038(w_010_038, w_001_002);
  and2 I010_040(w_010_040, w_003_089, w_002_017);
  or2  I010_041(w_010_041, w_007_091, w_008_309);
  nand2 I010_042(w_010_042, w_001_002, w_001_006);
  or2  I010_044(w_010_044, w_004_019, w_000_354);
  or2  I010_045(w_010_045, w_003_079, w_003_071);
  and2 I010_046(w_010_046, w_007_044, w_007_381);
  not1 I010_047(w_010_047, w_006_000);
  not1 I010_048(w_010_048, w_004_279);
  or2  I010_049(w_010_049, w_007_160, w_008_173);
  and2 I010_051(w_010_051, w_005_068, w_004_008);
  or2  I010_052(w_010_052, w_000_266, w_003_001);
  not1 I010_053(w_010_053, w_002_006);
  and2 I010_054(w_010_054, w_004_105, w_006_000);
  nand2 I010_055(w_010_055, w_001_001, w_002_008);
  nand2 I010_059(w_010_059, w_007_398, w_007_170);
  or2  I010_062(w_010_062, w_008_112, w_003_056);
  or2  I010_063(w_010_063, w_002_004, w_007_216);
  or2  I010_064(w_010_064, w_000_127, w_001_001);
  and2 I010_065(w_010_065, w_008_252, w_009_040);
  not1 I010_067(w_010_067, w_006_000);
  not1 I010_069(w_010_069, w_002_025);
  or2  I010_071(w_010_071, w_002_021, w_000_356);
  nand2 I010_072(w_010_072, w_005_049, w_001_000);
  or2  I010_073(w_010_073, w_009_112, w_007_080);
  or2  I010_075(w_010_075, w_001_003, w_001_004);
  nand2 I010_076(w_010_076, w_000_255, w_009_006);
  and2 I010_077(w_010_077, w_009_008, w_001_002);
  or2  I010_078(w_010_078, w_002_006, w_001_006);
  or2  I010_079(w_010_079, w_004_305, w_005_161);
  or2  I010_083(w_010_083, w_006_000, w_001_001);
  nand2 I010_087(w_010_087, w_009_173, w_006_000);
  not1 I010_089(w_010_089, w_009_034);
  and2 I010_094(w_010_094, w_007_121, w_008_254);
  or2  I010_096(w_010_096, w_000_358, w_003_019);
  and2 I010_097(w_010_097, w_001_002, w_009_038);
  or2  I010_098(w_010_098, w_004_438, w_003_023);
  nand2 I010_100(w_010_100, w_003_017, w_003_030);
  nand2 I010_101(w_010_101, w_002_012, w_008_223);
  and2 I010_103(w_010_103, w_008_031, w_004_142);
  or2  I010_104(w_010_104, w_003_010, w_004_249);
  or2  I010_107(w_010_107, w_000_359, w_004_054);
  nand2 I010_108(w_010_108, w_004_277, w_001_001);
  nand2 I010_112(w_010_112, w_008_067, w_004_354);
  or2  I010_115(w_010_115, w_005_022, w_002_018);
  or2  I010_116(w_010_116, w_009_194, w_001_001);
  not1 I010_119(w_010_119, w_007_343);
  not1 I010_120(w_010_120, w_000_360);
  nand2 I010_121(w_010_121, w_004_312, w_007_006);
  or2  I010_123(w_010_123, w_005_105, w_002_011);
  and2 I010_127(w_010_127, w_003_040, w_000_297);
  and2 I010_128(w_010_128, w_009_061, w_009_153);
  not1 I010_131(w_010_131, w_000_363);
  or2  I010_132(w_010_132, w_000_053, w_005_056);
  or2  I010_134(w_010_134, w_002_025, w_009_016);
  not1 I010_135(w_010_135, w_008_145);
  and2 I010_136(w_010_136, w_000_041, w_006_000);
  nand2 I010_137(w_010_137, w_003_009, w_005_211);
  nand2 I010_142(w_010_142, w_001_005, w_009_017);
  nand2 I010_144(w_010_144, w_001_005, w_003_052);
  not1 I010_145(w_010_145, w_006_000);
  nand2 I010_146(w_010_146, w_007_233, w_006_000);
  nand2 I010_150(w_010_150, w_000_164, w_005_060);
  nand2 I010_151(w_010_151, w_000_023, w_000_336);
  not1 I010_152(w_010_152, w_003_067);
  nand2 I010_153(w_010_153, w_009_047, w_008_062);
  or2  I010_158(w_010_158, w_002_015, w_007_285);
  not1 I010_159(w_010_159, w_006_000);
  and2 I010_162(w_010_162, w_006_000, w_008_008);
  or2  I010_163(w_010_163, w_000_292, w_003_076);
  not1 I010_170(w_010_170, w_007_092);
  or2  I010_172(w_010_172, w_004_010, w_005_017);
  or2  I010_174(w_010_174, w_009_007, w_002_011);
  and2 I010_175(w_010_175, w_009_168, w_007_355);
  or2  I010_176(w_010_176, w_001_005, w_009_198);
  and2 I010_178(w_010_178, w_007_297, w_001_002);
  not1 I010_179(w_010_179, w_007_092);
  or2  I010_180(w_010_180, w_007_371, w_002_000);
  and2 I010_181(w_010_181, w_002_000, w_009_089);
  not1 I010_185(w_010_185, w_000_236);
  nand2 I010_187(w_010_187, w_004_308, w_005_177);
  or2  I010_188(w_010_188, w_009_222, w_005_215);
  nand2 I010_189(w_010_189, w_006_000, w_001_003);
  not1 I010_190(w_010_190, w_009_090);
  nand2 I010_191(w_010_191, w_001_000, w_002_009);
  or2  I010_192(w_010_192, w_000_032, w_000_365);
  not1 I010_193(w_010_193, w_007_227);
  not1 I010_196(w_010_196, w_002_011);
  not1 I010_197(w_010_197, w_006_000);
  or2  I010_198(w_010_198, w_005_023, w_006_000);
  or2  I010_201(w_010_201, w_002_013, w_009_135);
  not1 I010_204(w_010_204, w_008_047);
  and2 I010_207(w_010_207, w_005_071, w_002_011);
  not1 I010_208(w_010_208, w_001_006);
  not1 I010_211(w_010_211, w_008_199);
  and2 I010_213(w_010_213, w_006_000, w_000_344);
  or2  I010_214(w_010_214, w_006_000, w_003_087);
  not1 I010_216(w_010_216, w_008_008);
  or2  I010_217(w_010_217, w_008_099, w_000_124);
  or2  I010_218(w_010_218, w_000_030, w_006_000);
  and2 I010_219(w_010_219, w_002_019, w_007_005);
  and2 I010_220(w_010_220, w_006_000, w_002_014);
  or2  I010_223(w_010_223, w_005_098, w_008_029);
  not1 I010_224(w_010_224, w_006_000);
  and2 I010_225(w_010_225, w_002_019, w_000_366);
  not1 I010_226(w_010_226, w_000_367);
  and2 I010_234(w_010_234, w_009_234, w_000_368);
  or2  I010_235(w_010_235, w_006_000, w_001_002);
  nand2 I010_236(w_010_236, w_002_026, w_004_259);
  and2 I010_240(w_010_240, w_005_005, w_007_315);
  or2  I010_241(w_010_241, w_008_161, w_004_141);
  not1 I010_244(w_010_244, w_002_021);
  not1 I010_246(w_010_246, w_007_051);
  nand2 I010_247(w_010_247, w_002_021, w_002_027);
  nand2 I010_251(w_010_251, w_000_204, w_009_177);
  nand2 I010_253(w_010_253, w_007_254, w_002_010);
  nand2 I010_254(w_010_254, w_004_141, w_008_177);
  not1 I010_255(w_010_255, w_005_088);
  or2  I010_256(w_010_256, w_006_000, w_002_008);
  not1 I010_258(w_010_258, w_002_016);
  or2  I010_260(w_010_260, w_007_138, w_003_071);
  or2  I010_261(w_010_261, w_000_213, w_002_003);
  nand2 I010_262(w_010_262, w_007_023, w_000_193);
  and2 I010_263(w_010_263, w_002_026, w_003_080);
  and2 I010_264(w_010_264, w_004_061, w_009_048);
  not1 I010_265(w_010_265, w_009_229);
  nand2 I010_266(w_010_266, w_001_001, w_008_120);
  nand2 I010_267(w_010_267, w_004_192, w_007_214);
  or2  I010_268(w_010_268, w_009_063, w_002_000);
  and2 I010_270(w_010_270, w_005_232, w_000_271);
  not1 I010_273(w_010_273, w_008_342);
  and2 I010_276(w_010_276, w_009_012, w_004_038);
  not1 I010_278(w_010_278, w_002_014);
  nand2 I010_281(w_010_281, w_000_371, w_005_106);
  nand2 I010_282(w_010_282, w_004_397, w_007_020);
  and2 I010_283(w_010_283, w_003_034, w_005_100);
  and2 I010_284(w_010_284, w_004_243, w_003_037);
  not1 I010_286(w_010_286, w_008_045);
  and2 I010_287(w_010_287, w_004_199, w_005_186);
  and2 I010_288(w_010_288, w_003_088, w_005_044);
  or2  I010_289(w_010_289, w_002_018, w_005_197);
  and2 I010_290(w_010_290, w_000_372, w_004_214);
  or2  I010_291(w_010_291, w_009_104, w_001_005);
  nand2 I010_292(w_010_292, w_006_000, w_003_046);
  or2  I010_294(w_010_294, w_005_106, w_001_000);
  and2 I010_298(w_010_298, w_000_091, w_001_002);
  not1 I010_303(w_010_303, w_008_149);
  not1 I010_304(w_010_304, w_009_232);
  not1 I010_306(w_010_306, w_001_005);
  and2 I010_307(w_010_307, w_004_233, w_009_186);
  and2 I010_309(w_010_309, w_002_011, w_000_373);
  nand2 I010_311(w_010_311, w_000_221, w_006_000);
  not1 I010_315(w_010_315, w_007_099);
  not1 I010_316(w_010_316, w_009_013);
  not1 I010_317(w_010_317, w_004_052);
  or2  I010_318(w_010_318, w_002_027, w_008_219);
  not1 I010_321(w_010_321, w_004_372);
  not1 I010_322(w_010_322, w_000_121);
  and2 I010_323(w_010_323, w_000_374, w_008_091);
  nand2 I010_325(w_010_325, w_008_258, w_009_128);
  nand2 I010_326(w_010_326, w_000_086, w_004_014);
  not1 I010_327(w_010_327, w_002_008);
  not1 I010_328(w_010_328, w_000_171);
  or2  I010_332(w_010_332, w_007_244, w_004_028);
  or2  I010_333(w_010_333, w_004_024, w_001_005);
  nand2 I010_334(w_010_334, w_007_281, w_000_001);
  not1 I010_336(w_010_336, w_000_194);
  not1 I010_337(w_010_337, w_005_223);
  and2 I010_338(w_010_338, w_009_014, w_009_031);
  nand2 I010_342(w_010_342, w_001_000, w_000_375);
  not1 I010_343(w_010_343, w_006_000);
  not1 I010_344(w_010_344, w_001_002);
  and2 I010_345(w_010_345, w_004_398, w_003_036);
  nand2 I010_346(w_010_346, w_003_066, w_004_447);
  nand2 I010_347(w_010_347, w_008_014, w_005_192);
  not1 I010_348(w_010_348, w_001_004);
  and2 I010_349(w_010_349, w_008_292, w_009_227);
  not1 I010_351(w_010_351, w_002_020);
  not1 I010_353(w_010_353, w_008_047);
  nand2 I010_354(w_010_354, w_004_130, w_000_306);
  not1 I010_357(w_010_357, w_002_026);
  or2  I010_359(w_010_359, w_002_019, w_003_093);
  not1 I010_361(w_010_361, w_006_000);
  and2 I010_362(w_010_362, w_002_024, w_009_108);
  or2  I010_364(w_010_364, w_009_047, w_005_152);
  nand2 I010_368(w_010_368, w_000_266, w_006_000);
  and2 I010_372(w_010_372, w_002_023, w_000_376);
  or2  I010_377(w_010_377, w_006_000, w_003_030);
  nand2 I010_379(w_010_379, w_000_377, w_008_062);
  or2  I010_380(w_010_380, w_008_003, w_009_079);
  and2 I010_381(w_010_381, w_000_228, w_000_378);
  nand2 I010_382(w_010_382, w_001_003, w_001_001);
  not1 I010_384(w_010_384, w_003_025);
  and2 I010_385(w_010_385, w_003_082, w_001_004);
  not1 I010_389(w_010_389, w_008_292);
  not1 I010_391(w_010_391, w_000_014);
  not1 I010_392(w_010_392, w_004_198);
  not1 I010_398(w_010_398, w_009_231);
  not1 I010_400(w_010_400, w_007_328);
  and2 I010_402(w_010_402, w_002_010, w_003_090);
  not1 I010_404(w_010_404, w_008_238);
  or2  I010_406(w_010_406, w_005_168, w_008_200);
  and2 I010_408(w_010_408, w_003_059, w_000_197);
  nand2 I010_410(w_010_410, w_008_005, w_001_005);
  and2 I010_412(w_010_412, w_004_224, w_006_000);
  or2  I010_413(w_010_413, w_005_081, w_003_037);
  not1 I010_416(w_010_416, w_003_039);
  or2  I010_417(w_010_417, w_001_002, w_005_144);
  and2 I010_418(w_010_418, w_003_100, w_001_003);
  or2  I010_422(w_010_422, w_005_067, w_002_017);
  not1 I010_423(w_010_423, w_005_101);
  not1 I010_425(w_010_425, w_002_006);
  or2  I010_427(w_010_427, w_005_108, w_000_381);
  not1 I010_429(w_010_429, w_003_095);
  and2 I010_431(w_010_431, w_004_289, w_009_144);
  nand2 I010_433(w_010_433, w_005_036, w_000_290);
  or2  I010_435(w_010_435, w_008_185, w_004_336);
  and2 I010_436(w_010_436, w_009_012, w_002_004);
  nand2 I010_438(w_010_438, w_005_032, w_009_003);
  and2 I010_441(w_010_441, w_002_020, w_005_058);
  nand2 I010_443(w_010_443, w_006_000, w_003_032);
  and2 I010_445(w_010_445, w_001_001, w_000_009);
  and2 I010_446(w_010_446, w_006_000, w_003_053);
  and2 I010_448(w_010_448, w_006_000, w_004_120);
  and2 I010_449(w_010_449, w_007_006, w_009_160);
  not1 I010_450(w_010_450, w_007_104);
  nand2 I010_451(w_010_451, w_008_128, w_006_000);
  nand2 I011_000(w_011_000, w_001_001, w_004_066);
  and2 I011_001(w_011_001, w_001_002, w_000_174);
  not1 I011_004(w_011_004, w_010_033);
  or2  I011_009(w_011_009, w_004_303, w_004_399);
  nand2 I011_011(w_011_011, w_006_000, w_002_017);
  or2  I011_012(w_011_012, w_001_003, w_009_144);
  and2 I011_014(w_011_014, w_005_175, w_009_031);
  not1 I011_015(w_011_015, w_007_190);
  or2  I011_016(w_011_016, w_010_089, w_007_071);
  not1 I011_017(w_011_017, w_003_057);
  or2  I011_018(w_011_018, w_009_046, w_003_068);
  or2  I011_019(w_011_019, w_004_386, w_007_381);
  or2  I011_020(w_011_020, w_001_002, w_008_079);
  and2 I011_021(w_011_021, w_000_254, w_006_000);
  and2 I011_022(w_011_022, w_000_382, w_001_002);
  or2  I011_023(w_011_023, w_006_000, w_002_008);
  not1 I011_025(w_011_025, w_005_163);
  nand2 I011_026(w_011_026, w_010_049, w_001_001);
  nand2 I011_027(w_011_027, w_000_115, w_003_049);
  and2 I011_028(w_011_028, w_001_006, w_007_226);
  nand2 I011_030(w_011_030, w_004_115, w_005_143);
  or2  I011_031(w_011_031, w_008_089, w_009_099);
  or2  I011_033(w_011_033, w_002_004, w_009_093);
  nand2 I011_034(w_011_034, w_008_292, w_006_000);
  not1 I011_035(w_011_035, w_003_005);
  or2  I011_036(w_011_036, w_001_004, w_002_006);
  or2  I011_037(w_011_037, w_008_034, w_010_298);
  not1 I011_038(w_011_038, w_006_000);
  or2  I011_039(w_011_039, w_009_153, w_000_145);
  and2 I011_041(w_011_041, w_000_264, w_001_006);
  nand2 I011_042(w_011_042, w_004_320, w_008_304);
  not1 I011_043(w_011_043, w_010_443);
  nand2 I011_045(w_011_045, w_002_019, w_009_237);
  not1 I011_047(w_011_047, w_009_044);
  nand2 I011_051(w_011_051, w_002_014, w_008_233);
  or2  I011_052(w_011_052, w_003_033, w_008_111);
  or2  I011_053(w_011_053, w_005_176, w_003_050);
  nand2 I011_054(w_011_054, w_001_001, w_009_088);
  not1 I011_055(w_011_055, w_004_458);
  or2  I011_056(w_011_056, w_002_021, w_001_004);
  and2 I011_057(w_011_057, w_007_041, w_010_291);
  and2 I011_058(w_011_058, w_005_024, w_002_019);
  or2  I011_059(w_011_059, w_008_130, w_000_021);
  and2 I011_060(w_011_060, w_003_025, w_006_000);
  nand2 I011_061(w_011_061, w_004_179, w_002_015);
  nand2 I011_063(w_011_063, w_006_000, w_009_129);
  nand2 I011_064(w_011_064, w_003_010, w_008_146);
  nand2 I011_066(w_011_066, w_001_005, w_002_001);
  nand2 I011_067(w_011_067, w_006_000, w_009_014);
  or2  I011_068(w_011_068, w_000_293, w_003_061);
  not1 I011_069(w_011_069, w_008_067);
  or2  I011_071(w_011_071, w_008_161, w_005_033);
  and2 I011_072(w_011_072, w_007_320, w_002_006);
  nand2 I011_073(w_011_073, w_004_372, w_002_024);
  and2 I011_076(w_011_076, w_003_071, w_006_000);
  and2 I011_077(w_011_077, w_002_015, w_001_002);
  or2  I011_078(w_011_078, w_008_043, w_003_034);
  or2  I011_079(w_011_079, w_003_031, w_010_425);
  or2  I011_080(w_011_080, w_005_150, w_010_220);
  nand2 I011_081(w_011_081, w_002_014, w_000_237);
  not1 I011_082(w_011_082, w_007_298);
  or2  I011_083(w_011_083, w_002_006, w_007_089);
  or2  I011_084(w_011_084, w_008_203, w_005_195);
  not1 I011_085(w_011_085, w_008_143);
  and2 I011_086(w_011_086, w_000_123, w_006_000);
  and2 I011_087(w_011_087, w_009_031, w_008_114);
  not1 I011_088(w_011_088, w_008_327);
  and2 I011_089(w_011_089, w_003_095, w_000_096);
  not1 I011_090(w_011_090, w_000_178);
  nand2 I011_091(w_011_091, w_000_331, w_004_183);
  or2  I011_092(w_011_092, w_005_029, w_009_025);
  not1 I011_093(w_011_093, w_009_000);
  or2  I011_095(w_011_095, w_002_004, w_010_075);
  and2 I011_096(w_011_096, w_002_020, w_001_003);
  not1 I011_097(w_011_097, w_010_181);
  or2  I011_098(w_011_098, w_000_012, w_009_103);
  or2  I011_099(w_011_099, w_003_021, w_004_312);
  or2  I011_100(w_011_100, w_000_164, w_002_019);
  or2  I011_101(w_011_101, w_001_001, w_005_241);
  not1 I011_102(w_011_102, w_004_421);
  or2  I011_104(w_011_104, w_007_180, w_000_005);
  and2 I011_106(w_011_106, w_007_075, w_008_297);
  and2 I011_108(w_011_108, w_003_051, w_005_193);
  nand2 I011_110(w_011_110, w_007_019, w_008_075);
  and2 I011_111(w_011_111, w_006_000, w_002_003);
  or2  I011_112(w_011_112, w_006_000, w_009_111);
  not1 I011_113(w_011_113, w_005_084);
  or2  I011_114(w_011_114, w_002_000, w_000_383);
  or2  I011_115(w_011_115, w_005_190, w_004_456);
  nand2 I011_116(w_011_116, w_007_225, w_008_085);
  or2  I011_117(w_011_117, w_003_001, w_000_316);
  nand2 I011_120(w_011_120, w_005_146, w_009_134);
  not1 I011_121(w_011_121, w_001_003);
  and2 I011_123(w_011_123, w_010_059, w_000_111);
  and2 I011_124(w_011_124, w_009_190, w_007_165);
  nand2 I011_125(w_011_125, w_000_030, w_005_189);
  or2  I011_126(w_011_126, w_001_004, w_007_363);
  nand2 I011_127(w_011_127, w_003_044, w_002_009);
  and2 I011_128(w_011_128, w_002_006, w_005_085);
  or2  I011_130(w_011_130, w_010_034, w_004_007);
  not1 I011_131(w_011_131, w_009_147);
  not1 I011_132(w_011_132, w_009_029);
  not1 I011_133(w_011_133, w_000_384);
  or2  I011_134(w_011_134, w_002_024, w_004_345);
  and2 I011_135(w_011_135, w_010_179, w_007_030);
  or2  I011_136(w_011_136, w_007_134, w_005_118);
  or2  I011_137(w_011_137, w_007_275, w_009_136);
  not1 I011_140(w_011_140, w_002_005);
  not1 I011_141(w_011_141, w_005_146);
  nand2 I011_142(w_011_142, w_004_078, w_009_021);
  nand2 I011_143(w_011_143, w_003_007, w_008_254);
  and2 I011_144(w_011_144, w_003_075, w_004_087);
  not1 I011_146(w_011_146, w_008_070);
  nand2 I011_150(w_011_150, w_009_045, w_003_061);
  nand2 I011_151(w_011_151, w_007_250, w_004_066);
  nand2 I011_152(w_011_152, w_000_386, w_010_236);
  not1 I011_153(w_011_153, w_001_004);
  or2  I011_155(w_011_155, w_009_144, w_003_066);
  and2 I011_156(w_011_156, w_003_061, w_009_027);
  and2 I011_159(w_011_159, w_000_170, w_005_007);
  nand2 I011_160(w_011_160, w_003_067, w_006_000);
  nand2 I011_161(w_011_161, w_001_006, w_003_088);
  nand2 I011_163(w_011_163, w_002_013, w_002_016);
  nand2 I011_164(w_011_164, w_009_092, w_006_000);
  not1 I011_166(w_011_166, w_003_051);
  not1 I011_169(w_011_169, w_008_152);
  or2  I011_177(w_011_177, w_010_398, w_009_002);
  or2  I011_178(w_011_178, w_002_000, w_000_293);
  or2  I011_179(w_011_179, w_008_039, w_009_049);
  not1 I011_181(w_011_181, w_001_000);
  nand2 I011_182(w_011_182, w_000_112, w_001_002);
  nand2 I011_183(w_011_183, w_007_329, w_007_163);
  nand2 I011_186(w_011_186, w_005_226, w_008_161);
  and2 I011_187(w_011_187, w_002_023, w_004_311);
  or2  I011_188(w_011_188, w_003_077, w_003_025);
  or2  I011_189(w_011_189, w_003_053, w_005_038);
  or2  I011_192(w_011_192, w_003_087, w_004_386);
  and2 I011_194(w_011_194, w_000_224, w_002_018);
  and2 I011_196(w_011_196, w_004_394, w_001_000);
  not1 I011_197(w_011_197, w_005_107);
  not1 I011_200(w_011_200, w_001_005);
  nand2 I011_201(w_011_201, w_006_000, w_009_178);
  and2 I011_204(w_011_204, w_006_000, w_000_075);
  and2 I011_205(w_011_205, w_007_253, w_000_128);
  not1 I011_206(w_011_206, w_009_021);
  or2  I011_207(w_011_207, w_008_041, w_008_331);
  and2 I011_211(w_011_211, w_002_013, w_007_120);
  or2  I011_213(w_011_213, w_003_097, w_008_342);
  or2  I011_214(w_011_214, w_003_026, w_000_279);
  or2  I011_215(w_011_215, w_003_015, w_009_185);
  nand2 I011_218(w_011_218, w_010_007, w_010_021);
  not1 I011_219(w_011_219, w_004_426);
  nand2 I011_220(w_011_220, w_006_000, w_009_073);
  or2  I011_221(w_011_221, w_010_451, w_006_000);
  or2  I011_222(w_011_222, w_010_045, w_010_402);
  or2  I011_224(w_011_224, w_004_006, w_004_010);
  and2 I011_226(w_011_226, w_005_238, w_007_075);
  nand2 I011_228(w_011_228, w_003_044, w_008_199);
  and2 I011_230(w_011_230, w_004_410, w_008_324);
  nand2 I011_231(w_011_231, w_002_014, w_006_000);
  and2 I011_232(w_011_232, w_005_133, w_000_187);
  and2 I011_233(w_011_233, w_007_115, w_004_274);
  and2 I011_234(w_011_234, w_006_000, w_001_004);
  or2  I011_238(w_011_238, w_009_221, w_004_020);
  nand2 I011_242(w_011_242, w_003_064, w_009_125);
  and2 I011_246(w_011_246, w_003_014, w_010_346);
  nand2 I011_249(w_011_249, w_008_255, w_006_000);
  or2  I011_251(w_011_251, w_001_006, w_006_000);
  or2  I011_253(w_011_253, w_002_018, w_005_145);
  not1 I011_254(w_011_254, w_006_000);
  not1 I011_257(w_011_257, w_005_109);
  or2  I011_268(w_011_268, w_006_000, w_000_307);
  and2 I011_269(w_011_269, w_005_163, w_009_106);
  not1 I011_272(w_011_272, w_004_025);
  not1 I011_273(w_011_273, w_001_003);
  nand2 I011_276(w_011_276, w_004_305, w_007_031);
  and2 I011_278(w_011_278, w_000_246, w_008_168);
  or2  I011_279(w_011_279, w_007_306, w_010_266);
  or2  I011_280(w_011_280, w_000_268, w_000_389);
  nand2 I011_282(w_011_282, w_008_329, w_004_130);
  and2 I011_284(w_011_284, w_009_064, w_009_144);
  and2 I011_285(w_011_285, w_004_050, w_001_001);
  and2 I011_286(w_011_286, w_001_001, w_008_253);
  or2  I011_287(w_011_287, w_006_000, w_003_004);
  or2  I011_289(w_011_289, w_001_004, w_003_074);
  not1 I011_291(w_011_291, w_008_269);
  and2 I011_292(w_011_292, w_008_001, w_000_032);
  and2 I011_294(w_011_294, w_010_016, w_000_045);
  or2  I011_295(w_011_295, w_008_150, w_007_377);
  or2  I011_296(w_011_296, w_000_304, w_003_073);
  and2 I011_297(w_011_297, w_005_061, w_004_225);
  not1 I011_300(w_011_300, w_002_004);
  not1 I011_301(w_011_301, w_002_001);
  and2 I011_303(w_011_303, w_005_101, w_007_213);
  nand2 I011_304(w_011_304, w_007_341, w_004_273);
  not1 I011_308(w_011_308, w_003_052);
  nand2 I011_309(w_011_309, w_000_017, w_005_196);
  and2 I011_312(w_011_312, w_004_452, w_001_003);
  not1 I011_315(w_011_315, w_000_033);
  and2 I011_317(w_011_317, w_009_108, w_006_000);
  nand2 I011_318(w_011_318, w_004_132, w_009_046);
  or2  I011_319(w_011_319, w_008_034, w_001_000);
  nand2 I011_320(w_011_320, w_009_128, w_005_224);
  and2 I011_321(w_011_321, w_007_243, w_009_121);
  or2  I011_323(w_011_323, w_005_162, w_001_006);
  or2  I011_327(w_011_327, w_005_077, w_010_244);
  not1 I011_329(w_011_329, w_008_150);
  nand2 I011_331(w_011_331, w_008_080, w_000_123);
  not1 I011_332(w_011_332, w_008_098);
  not1 I011_333(w_011_333, w_003_027);
  not1 I011_334(w_011_334, w_007_026);
  nand2 I011_335(w_011_335, w_008_175, w_004_255);
  not1 I011_336(w_011_336, w_000_390);
  not1 I011_337(w_011_337, w_009_236);
  and2 I011_339(w_011_339, w_006_000, w_003_039);
  or2  I011_340(w_011_340, w_009_094, w_008_073);
  not1 I011_342(w_011_342, w_007_377);
  nand2 I012_000(w_012_000, w_011_111, w_008_027);
  and2 I012_001(w_012_001, w_010_449, w_010_158);
  not1 I012_002(w_012_002, w_002_023);
  not1 I012_003(w_012_003, w_000_323);
  or2  I012_004(w_012_004, w_006_000, w_011_142);
  nand2 I012_005(w_012_005, w_003_004, w_006_000);
  and2 I012_006(w_012_006, w_004_113, w_002_015);
  and2 I012_007(w_012_007, w_001_004, w_000_063);
  and2 I012_010(w_012_010, w_007_087, w_001_003);
  or2  I012_012(w_012_012, w_008_070, w_003_069);
  or2  I012_013(w_012_013, w_007_035, w_003_050);
  nand2 I012_014(w_012_014, w_008_012, w_000_219);
  not1 I012_015(w_012_015, w_003_028);
  not1 I012_016(w_012_016, w_004_194);
  and2 I012_017(w_012_017, w_001_003, w_003_083);
  and2 I012_018(w_012_018, w_008_239, w_005_230);
  and2 I012_019(w_012_019, w_001_000, w_003_001);
  and2 I012_020(w_012_020, w_010_342, w_007_048);
  or2  I012_021(w_012_021, w_008_317, w_001_004);
  not1 I012_023(w_012_023, w_001_003);
  or2  I012_024(w_012_024, w_005_103, w_001_003);
  not1 I012_025(w_012_025, w_007_196);
  not1 I012_026(w_012_026, w_000_391);
  or2  I012_027(w_012_027, w_003_026, w_007_373);
  and2 I012_028(w_012_028, w_004_343, w_004_225);
  and2 I012_029(w_012_029, w_003_020, w_001_001);
  or2  I012_030(w_012_030, w_010_273, w_007_200);
  not1 I012_031(w_012_031, w_004_303);
  nand2 I012_032(w_012_032, w_001_000, w_002_014);
  not1 I012_034(w_012_034, w_011_004);
  not1 I012_035(w_012_035, w_008_199);
  not1 I012_036(w_012_036, w_005_006);
  or2  I012_038(w_012_038, w_007_154, w_006_000);
  not1 I012_039(w_012_039, w_000_370);
  or2  I012_040(w_012_040, w_003_022, w_002_014);
  not1 I012_041(w_012_041, w_005_112);
  and2 I012_042(w_012_042, w_009_143, w_006_000);
  nand2 I012_043(w_012_043, w_001_005, w_006_000);
  and2 I012_045(w_012_045, w_002_006, w_000_189);
  and2 I012_046(w_012_046, w_006_000, w_004_465);
  nand2 I012_048(w_012_048, w_009_147, w_003_058);
  not1 I012_049(w_012_049, w_001_004);
  not1 I012_050(w_012_050, w_002_020);
  nand2 I012_052(w_012_052, w_005_006, w_007_025);
  not1 I012_053(w_012_053, w_002_009);
  nand2 I012_054(w_012_054, w_011_286, w_007_092);
  not1 I012_055(w_012_055, w_005_170);
  nand2 I012_056(w_012_056, w_000_392, w_009_008);
  nand2 I012_057(w_012_057, w_009_002, w_006_000);
  and2 I012_060(w_012_060, w_001_002, w_003_024);
  not1 I012_061(w_012_061, w_010_116);
  or2  I012_063(w_012_063, w_005_121, w_009_196);
  nand2 I012_065(w_012_065, w_007_172, w_006_000);
  and2 I012_067(w_012_067, w_009_155, w_003_077);
  and2 I012_068(w_012_068, w_005_145, w_000_188);
  and2 I012_070(w_012_070, w_004_367, w_006_000);
  not1 I012_071(w_012_071, w_009_226);
  not1 I012_073(w_012_073, w_003_070);
  not1 I012_074(w_012_074, w_000_284);
  not1 I012_077(w_012_077, w_003_043);
  and2 I012_080(w_012_080, w_007_352, w_000_038);
  nand2 I012_081(w_012_081, w_001_001, w_003_085);
  or2  I012_083(w_012_083, w_006_000, w_004_029);
  or2  I012_084(w_012_084, w_004_325, w_000_393);
  nand2 I012_086(w_012_086, w_000_354, w_009_229);
  and2 I012_088(w_012_088, w_006_000, w_003_093);
  or2  I012_089(w_012_089, w_009_021, w_007_270);
  nand2 I012_090(w_012_090, w_008_126, w_008_236);
  and2 I012_091(w_012_091, w_008_282, w_000_176);
  and2 I012_092(w_012_092, w_007_104, w_007_055);
  or2  I012_094(w_012_094, w_010_289, w_008_109);
  or2  I012_096(w_012_096, w_009_010, w_003_092);
  not1 I012_097(w_012_097, w_007_350);
  or2  I012_098(w_012_098, w_007_027, w_005_146);
  nand2 I012_099(w_012_099, w_004_106, w_011_211);
  and2 I012_101(w_012_101, w_009_146, w_009_021);
  not1 I012_103(w_012_103, w_003_089);
  nand2 I012_108(w_012_108, w_002_019, w_011_186);
  and2 I012_109(w_012_109, w_011_183, w_002_023);
  not1 I012_110(w_012_110, w_007_138);
  and2 I012_113(w_012_113, w_000_394, w_001_000);
  not1 I012_114(w_012_114, w_007_035);
  nand2 I012_116(w_012_116, w_000_030, w_010_046);
  or2  I012_119(w_012_119, w_004_155, w_001_002);
  nand2 I012_122(w_012_122, w_002_010, w_002_002);
  nand2 I012_125(w_012_125, w_005_124, w_006_000);
  not1 I012_126(w_012_126, w_010_028);
  nand2 I012_127(w_012_127, w_006_000, w_005_169);
  nand2 I012_131(w_012_131, w_009_113, w_004_286);
  not1 I012_132(w_012_132, w_010_015);
  or2  I012_133(w_012_133, w_011_201, w_007_276);
  or2  I012_135(w_012_135, w_001_002, w_001_003);
  and2 I012_138(w_012_138, w_002_003, w_000_388);
  nand2 I012_143(w_012_143, w_008_208, w_000_395);
  and2 I012_144(w_012_144, w_008_191, w_011_089);
  or2  I012_146(w_012_146, w_001_002, w_003_093);
  or2  I012_147(w_012_147, w_004_031, w_005_113);
  or2  I012_149(w_012_149, w_003_077, w_002_020);
  or2  I012_151(w_012_151, w_010_135, w_001_001);
  not1 I012_158(w_012_158, w_011_079);
  or2  I012_159(w_012_159, w_006_000, w_001_000);
  and2 I012_160(w_012_160, w_006_000, w_009_185);
  or2  I012_161(w_012_161, w_002_019, w_001_001);
  and2 I012_165(w_012_165, w_003_009, w_009_203);
  nand2 I012_166(w_012_166, w_002_021, w_007_052);
  not1 I012_169(w_012_169, w_011_337);
  or2  I012_170(w_012_170, w_008_209, w_000_039);
  not1 I012_171(w_012_171, w_010_004);
  or2  I012_174(w_012_174, w_010_281, w_009_175);
  not1 I012_175(w_012_175, w_008_307);
  nand2 I012_176(w_012_176, w_001_006, w_007_242);
  not1 I012_177(w_012_177, w_003_099);
  nand2 I012_178(w_012_178, w_006_000, w_001_003);
  and2 I012_180(w_012_180, w_005_161, w_005_151);
  not1 I012_181(w_012_181, w_008_087);
  nand2 I012_182(w_012_182, w_009_155, w_007_248);
  or2  I012_184(w_012_184, w_007_263, w_001_005);
  nand2 I012_186(w_012_186, w_007_135, w_001_001);
  nand2 I012_187(w_012_187, w_008_104, w_004_213);
  nand2 I012_189(w_012_189, w_006_000, w_010_078);
  nand2 I012_191(w_012_191, w_007_026, w_008_166);
  and2 I012_195(w_012_195, w_008_047, w_010_449);
  or2  I012_197(w_012_197, w_011_111, w_004_426);
  not1 I012_200(w_012_200, w_004_168);
  or2  I012_201(w_012_201, w_006_000, w_000_283);
  or2  I012_205(w_012_205, w_008_080, w_004_011);
  and2 I012_211(w_012_211, w_006_000, w_002_013);
  nand2 I012_212(w_012_212, w_010_253, w_007_357);
  or2  I012_214(w_012_214, w_007_040, w_006_000);
  and2 I012_215(w_012_215, w_004_128, w_011_221);
  and2 I012_217(w_012_217, w_010_213, w_000_220);
  not1 I012_218(w_012_218, w_006_000);
  or2  I012_219(w_012_219, w_005_147, w_004_094);
  and2 I012_220(w_012_220, w_009_050, w_010_246);
  or2  I012_221(w_012_221, w_005_191, w_008_045);
  nand2 I012_222(w_012_222, w_004_019, w_006_000);
  or2  I012_223(w_012_223, w_001_002, w_009_183);
  and2 I012_225(w_012_225, w_004_469, w_003_076);
  nand2 I012_226(w_012_226, w_011_146, w_007_285);
  nand2 I012_227(w_012_227, w_001_005, w_011_337);
  or2  I012_230(w_012_230, w_011_073, w_001_006);
  nand2 I012_234(w_012_234, w_004_312, w_001_001);
  or2  I012_236(w_012_236, w_004_046, w_002_025);
  and2 I012_238(w_012_238, w_007_147, w_008_028);
  not1 I012_239(w_012_239, w_009_116);
  nand2 I012_241(w_012_241, w_008_157, w_004_345);
  and2 I012_245(w_012_245, w_009_091, w_004_383);
  or2  I012_248(w_012_248, w_010_284, w_005_139);
  and2 I012_249(w_012_249, w_004_032, w_002_015);
  not1 I012_250(w_012_250, w_007_015);
  and2 I012_253(w_012_253, w_011_238, w_007_086);
  not1 I012_255(w_012_255, w_000_397);
  nand2 I012_256(w_012_256, w_004_459, w_001_002);
  nand2 I012_258(w_012_258, w_007_089, w_000_247);
  and2 I012_260(w_012_260, w_007_143, w_005_156);
  not1 I012_261(w_012_261, w_000_344);
  and2 I012_262(w_012_262, w_004_271, w_003_038);
  not1 I012_263(w_012_263, w_005_048);
  nand2 I012_265(w_012_265, w_009_050, w_011_113);
  not1 I012_266(w_012_266, w_008_090);
  not1 I012_270(w_012_270, w_008_137);
  not1 I012_272(w_012_272, w_000_008);
  and2 I012_275(w_012_275, w_009_018, w_003_003);
  nand2 I012_277(w_012_277, w_000_398, w_010_145);
  not1 I012_278(w_012_278, w_003_090);
  or2  I012_279(w_012_279, w_003_053, w_004_130);
  nand2 I012_280(w_012_280, w_004_020, w_007_045);
  nand2 I012_282(w_012_282, w_005_189, w_010_260);
  or2  I012_283(w_012_283, w_004_378, w_001_005);
  or2  I012_284(w_012_284, w_002_018, w_004_219);
  and2 I012_285(w_012_285, w_011_014, w_009_132);
  or2  I012_286(w_012_286, w_002_001, w_004_410);
  and2 I012_290(w_012_290, w_009_222, w_001_003);
  not1 I012_291(w_012_291, w_005_026);
  not1 I012_293(w_012_293, w_010_348);
  not1 I012_294(w_012_294, w_008_048);
  or2  I012_295(w_012_295, w_004_167, w_005_005);
  or2  I012_296(w_012_296, w_007_030, w_001_002);
  not1 I012_298(w_012_298, w_000_248);
  and2 I012_300(w_012_300, w_007_210, w_002_019);
  nand2 I012_303(w_012_303, w_002_003, w_007_252);
  or2  I012_309(w_012_309, w_006_000, w_005_146);
  nand2 I012_310(w_012_310, w_007_005, w_001_002);
  not1 I012_312(w_012_312, w_001_005);
  or2  I012_313(w_012_313, w_001_000, w_002_016);
  or2  I012_314(w_012_314, w_010_290, w_000_030);
  or2  I012_315(w_012_315, w_006_000, w_003_011);
  and2 I012_318(w_012_318, w_003_090, w_006_000);
  and2 I012_320(w_012_320, w_004_086, w_005_119);
  and2 I012_321(w_012_321, w_009_001, w_005_178);
  or2  I012_322(w_012_322, w_008_146, w_004_370);
  nand2 I012_324(w_012_324, w_003_012, w_011_159);
  nand2 I012_325(w_012_325, w_006_000, w_009_196);
  not1 I012_326(w_012_326, w_001_001);
  or2  I012_328(w_012_328, w_006_000, w_005_066);
  and2 I012_330(w_012_330, w_006_000, w_003_035);
  not1 I012_333(w_012_333, w_001_000);
  or2  I012_336(w_012_336, w_008_300, w_001_001);
  not1 I012_337(w_012_337, w_005_136);
  not1 I012_339(w_012_339, w_006_000);
  nand2 I012_340(w_012_340, w_003_089, w_004_209);
  or2  I012_341(w_012_341, w_000_162, w_000_098);
  and2 I012_344(w_012_344, w_005_040, w_010_214);
  not1 I012_345(w_012_345, w_007_396);
  or2  I012_347(w_012_347, w_008_239, w_002_009);
  or2  I012_348(w_012_348, w_002_023, w_002_010);
  or2  I012_349(w_012_349, w_004_368, w_000_399);
  not1 I012_350(w_012_350, w_008_345);
  nand2 I012_353(w_012_353, w_004_132, w_004_417);
  nand2 I012_356(w_012_356, w_010_344, w_006_000);
  or2  I012_357(w_012_357, w_009_232, w_003_016);
  and2 I012_358(w_012_358, w_011_218, w_004_115);
  or2  I012_359(w_012_359, w_004_372, w_009_126);
  or2  I012_362(w_012_362, w_000_096, w_005_182);
  not1 I012_363(w_012_363, w_006_000);
  nand2 I012_364(w_012_364, w_009_059, w_007_356);
  nand2 I012_365(w_012_365, w_000_324, w_000_260);
  and2 I012_366(w_012_366, w_009_124, w_009_077);
  and2 I012_367(w_012_367, w_004_137, w_005_012);
  and2 I012_368(w_012_368, w_005_110, w_005_233);
  not1 I012_369(w_012_369, w_002_023);
  not1 I012_373(w_012_373, w_005_114);
  nand2 I012_374(w_012_374, w_002_027, w_007_360);
  and2 I012_379(w_012_379, w_005_092, w_008_030);
  nand2 I012_380(w_012_380, w_003_068, w_011_121);
  or2  I012_382(w_012_382, w_004_247, w_008_236);
  not1 I013_000(w_013_000, w_007_356);
  nand2 I013_001(w_013_001, w_002_020, w_008_032);
  and2 I013_005(w_013_005, w_001_004, w_003_075);
  or2  I013_006(w_013_006, w_009_170, w_001_001);
  not1 I013_007(w_013_007, w_008_321);
  or2  I013_008(w_013_008, w_000_085, w_009_158);
  and2 I013_009(w_013_009, w_005_231, w_001_004);
  or2  I013_010(w_013_010, w_010_307, w_004_339);
  and2 I013_011(w_013_011, w_004_295, w_000_223);
  nand2 I013_012(w_013_012, w_005_002, w_004_263);
  not1 I013_013(w_013_013, w_008_031);
  and2 I013_014(w_013_014, w_003_096, w_005_222);
  or2  I013_017(w_013_017, w_012_099, w_011_187);
  or2  I013_018(w_013_018, w_001_003, w_000_158);
  and2 I013_019(w_013_019, w_006_000, w_012_031);
  nand2 I013_020(w_013_020, w_003_041, w_011_041);
  not1 I013_022(w_013_022, w_006_000);
  not1 I013_023(w_013_023, w_009_000);
  nand2 I013_024(w_013_024, w_009_127, w_010_094);
  not1 I013_025(w_013_025, w_004_372);
  not1 I013_027(w_013_027, w_002_013);
  not1 I013_028(w_013_028, w_012_265);
  and2 I013_030(w_013_030, w_003_012, w_012_275);
  nand2 I013_032(w_013_032, w_001_004, w_003_014);
  nand2 I013_033(w_013_033, w_010_029, w_003_016);
  nand2 I013_034(w_013_034, w_005_000, w_010_071);
  not1 I013_035(w_013_035, w_001_006);
  and2 I013_036(w_013_036, w_005_242, w_003_101);
  and2 I013_037(w_013_037, w_002_023, w_011_295);
  or2  I013_038(w_013_038, w_008_037, w_002_011);
  or2  I013_039(w_013_039, w_007_203, w_008_130);
  and2 I013_040(w_013_040, w_000_401, w_008_245);
  nand2 I013_041(w_013_041, w_006_000, w_000_259);
  or2  I013_043(w_013_043, w_005_159, w_001_005);
  not1 I013_044(w_013_044, w_003_045);
  nand2 I013_046(w_013_046, w_003_063, w_008_282);
  nand2 I013_047(w_013_047, w_003_073, w_012_211);
  and2 I013_049(w_013_049, w_006_000, w_012_230);
  not1 I013_050(w_013_050, w_000_340);
  and2 I013_051(w_013_051, w_006_000, w_000_325);
  or2  I013_052(w_013_052, w_008_212, w_011_141);
  or2  I013_053(w_013_053, w_006_000, w_009_083);
  not1 I013_054(w_013_054, w_011_042);
  not1 I013_055(w_013_055, w_012_060);
  not1 I013_057(w_013_057, w_001_003);
  or2  I013_059(w_013_059, w_003_016, w_006_000);
  and2 I013_060(w_013_060, w_005_085, w_009_003);
  not1 I013_061(w_013_061, w_006_000);
  or2  I013_062(w_013_062, w_003_035, w_012_282);
  and2 I013_063(w_013_063, w_005_162, w_009_178);
  nand2 I013_065(w_013_065, w_002_005, w_001_002);
  not1 I013_066(w_013_066, w_008_075);
  not1 I013_068(w_013_068, w_000_107);
  or2  I013_071(w_013_071, w_003_088, w_003_016);
  and2 I013_073(w_013_073, w_009_001, w_012_127);
  nand2 I013_075(w_013_075, w_000_403, w_008_256);
  and2 I013_080(w_013_080, w_002_021, w_001_001);
  not1 I013_081(w_013_081, w_003_008);
  not1 I013_082(w_013_082, w_005_010);
  and2 I013_083(w_013_083, w_008_090, w_009_015);
  and2 I013_084(w_013_084, w_002_027, w_002_014);
  or2  I013_087(w_013_087, w_005_112, w_009_084);
  nand2 I013_088(w_013_088, w_001_000, w_000_315);
  or2  I013_089(w_013_089, w_005_231, w_002_021);
  and2 I013_090(w_013_090, w_003_088, w_010_423);
  not1 I013_091(w_013_091, w_002_015);
  nand2 I013_093(w_013_093, w_012_040, w_008_113);
  and2 I013_094(w_013_094, w_007_030, w_006_000);
  or2  I013_095(w_013_095, w_008_176, w_002_021);
  nand2 I013_096(w_013_096, w_006_000, w_004_219);
  nand2 I013_097(w_013_097, w_001_004, w_008_026);
  nand2 I013_099(w_013_099, w_007_276, w_000_254);
  or2  I013_100(w_013_100, w_001_005, w_008_321);
  or2  I013_101(w_013_101, w_001_002, w_012_285);
  nand2 I013_102(w_013_102, w_005_207, w_009_001);
  nand2 I013_103(w_013_103, w_010_247, w_001_003);
  and2 I013_104(w_013_104, w_001_005, w_012_212);
  nand2 I013_105(w_013_105, w_012_330, w_011_160);
  and2 I013_106(w_013_106, w_011_027, w_007_061);
  and2 I013_108(w_013_108, w_005_177, w_003_071);
  not1 I013_109(w_013_109, w_001_005);
  or2  I013_110(w_013_110, w_002_014, w_007_376);
  nand2 I013_112(w_013_112, w_012_349, w_007_189);
  not1 I013_113(w_013_113, w_004_406);
  nand2 I013_116(w_013_116, w_003_033, w_011_113);
  not1 I013_117(w_013_117, w_003_091);
  and2 I013_118(w_013_118, w_010_304, w_003_012);
  or2  I013_119(w_013_119, w_006_000, w_004_418);
  not1 I013_120(w_013_120, w_007_164);
  nand2 I013_122(w_013_122, w_011_025, w_004_439);
  and2 I013_123(w_013_123, w_008_324, w_001_006);
  not1 I013_124(w_013_124, w_006_000);
  nand2 I013_126(w_013_126, w_004_082, w_004_125);
  nand2 I013_127(w_013_127, w_003_083, w_009_024);
  or2  I013_129(w_013_129, w_003_035, w_004_328);
  or2  I013_132(w_013_132, w_004_030, w_007_090);
  and2 I013_133(w_013_133, w_000_120, w_012_286);
  and2 I013_134(w_013_134, w_008_162, w_005_037);
  and2 I013_135(w_013_135, w_010_353, w_005_136);
  not1 I013_140(w_013_140, w_008_128);
  or2  I013_141(w_013_141, w_011_045, w_007_014);
  nand2 I013_142(w_013_142, w_010_015, w_007_224);
  not1 I013_144(w_013_144, w_005_121);
  or2  I013_145(w_013_145, w_005_184, w_006_000);
  not1 I013_146(w_013_146, w_006_000);
  not1 I013_147(w_013_147, w_002_001);
  or2  I013_148(w_013_148, w_006_000, w_010_201);
  and2 I013_149(w_013_149, w_010_192, w_005_134);
  nand2 I013_150(w_013_150, w_011_073, w_011_031);
  or2  I013_151(w_013_151, w_006_000, w_003_044);
  not1 I013_152(w_013_152, w_008_089);
  and2 I013_153(w_013_153, w_005_029, w_006_000);
  and2 I013_154(w_013_154, w_008_180, w_007_359);
  not1 I013_155(w_013_155, w_004_060);
  not1 I013_158(w_013_158, w_012_054);
  not1 I013_159(w_013_159, w_004_071);
  and2 I013_160(w_013_160, w_009_164, w_010_343);
  and2 I013_161(w_013_161, w_003_000, w_001_006);
  nand2 I013_162(w_013_162, w_006_000, w_005_030);
  or2  I013_163(w_013_163, w_009_096, w_004_183);
  not1 I013_164(w_013_164, w_010_323);
  nand2 I013_165(w_013_165, w_005_180, w_005_153);
  and2 I013_166(w_013_166, w_010_224, w_002_026);
  and2 I013_167(w_013_167, w_001_004, w_001_000);
  or2  I013_168(w_013_168, w_004_023, w_001_002);
  not1 I013_169(w_013_169, w_007_049);
  and2 I013_171(w_013_171, w_008_038, w_000_404);
  not1 I013_172(w_013_172, w_008_077);
  not1 I013_173(w_013_173, w_007_147);
  not1 I013_174(w_013_174, w_002_016);
  nand2 I013_175(w_013_175, w_010_197, w_000_261);
  or2  I013_176(w_013_176, w_009_190, w_000_405);
  or2  I013_177(w_013_177, w_008_115, w_012_226);
  and2 I013_180(w_013_180, w_011_321, w_000_348);
  nand2 I013_181(w_013_181, w_002_004, w_001_001);
  or2  I013_182(w_013_182, w_003_013, w_003_052);
  nand2 I013_183(w_013_183, w_004_254, w_000_127);
  and2 I013_184(w_013_184, w_012_205, w_010_136);
  and2 I013_185(w_013_185, w_009_211, w_003_087);
  and2 I013_186(w_013_186, w_009_151, w_009_045);
  or2  I013_187(w_013_187, w_004_043, w_005_222);
  nand2 I013_188(w_013_188, w_008_098, w_009_011);
  not1 I013_189(w_013_189, w_005_201);
  or2  I013_190(w_013_190, w_007_328, w_009_172);
  not1 I013_191(w_013_191, w_006_000);
  not1 I013_192(w_013_192, w_004_109);
  and2 I013_193(w_013_193, w_003_041, w_002_003);
  not1 I013_194(w_013_194, w_011_068);
  not1 I013_195(w_013_195, w_011_098);
  or2  I013_196(w_013_196, w_012_029, w_000_187);
  or2  I013_197(w_013_197, w_000_255, w_001_002);
  or2  I013_199(w_013_199, w_004_395, w_001_006);
  nand2 I013_200(w_013_200, w_004_054, w_006_000);
  and2 I013_201(w_013_201, w_004_127, w_005_178);
  not1 I013_204(w_013_204, w_010_112);
  not1 I013_205(w_013_205, w_005_245);
  nand2 I013_207(w_013_207, w_005_034, w_002_020);
  nand2 I013_208(w_013_208, w_006_000, w_008_168);
  not1 I013_210(w_013_210, w_011_320);
  not1 I013_211(w_013_211, w_005_070);
  not1 I013_213(w_013_213, w_005_199);
  not1 I013_214(w_013_214, w_010_021);
  nand2 I013_215(w_013_215, w_007_076, w_003_052);
  nand2 I013_217(w_013_217, w_007_100, w_011_092);
  or2  I013_218(w_013_218, w_011_301, w_006_000);
  or2  I013_220(w_013_220, w_008_102, w_002_018);
  nand2 I013_221(w_013_221, w_003_094, w_011_037);
  not1 I013_222(w_013_222, w_001_000);
  or2  I013_223(w_013_223, w_006_000, w_012_053);
  nand2 I013_224(w_013_224, w_012_114, w_000_157);
  not1 I013_225(w_013_225, w_008_258);
  or2  I013_226(w_013_226, w_010_013, w_008_098);
  not1 I013_227(w_013_227, w_005_145);
  or2  I013_228(w_013_228, w_000_173, w_010_132);
  and2 I013_229(w_013_229, w_003_039, w_011_076);
  nand2 I013_231(w_013_231, w_012_032, w_012_280);
  not1 I013_232(w_013_232, w_009_152);
  not1 I013_235(w_013_235, w_008_270);
  nand2 I013_239(w_013_239, w_000_017, w_006_000);
  or2  I013_243(w_013_243, w_006_000, w_007_105);
  not1 I013_245(w_013_245, w_001_005);
  nand2 I013_246(w_013_246, w_007_070, w_011_086);
  nand2 I013_248(w_013_248, w_009_001, w_010_132);
  and2 I013_250(w_013_250, w_003_063, w_006_000);
  not1 I013_253(w_013_253, w_009_050);
  not1 I013_255(w_013_255, w_000_075);
  not1 I013_261(w_013_261, w_012_001);
  or2  I013_264(w_013_264, w_004_328, w_006_000);
  nand2 I013_265(w_013_265, w_000_408, w_000_409);
  nand2 I013_266(w_013_266, w_012_373, w_007_072);
  or2  I013_267(w_013_267, w_010_187, w_001_002);
  or2  I013_268(w_013_268, w_000_157, w_003_004);
  nand2 I014_001(w_014_001, w_013_218, w_011_207);
  nand2 I014_002(w_014_002, w_010_174, w_003_006);
  or2  I014_005(w_014_005, w_009_007, w_009_164);
  and2 I014_006(w_014_006, w_005_082, w_001_000);
  and2 I014_007(w_014_007, w_007_278, w_006_000);
  or2  I014_008(w_014_008, w_003_037, w_008_083);
  and2 I014_009(w_014_009, w_011_053, w_012_004);
  not1 I014_010(w_014_010, w_011_272);
  or2  I014_011(w_014_011, w_008_079, w_000_145);
  or2  I014_013(w_014_013, w_012_038, w_000_017);
  nand2 I014_014(w_014_014, w_004_199, w_005_078);
  nand2 I014_016(w_014_016, w_000_410, w_003_034);
  nand2 I014_017(w_014_017, w_006_000, w_010_144);
  and2 I014_018(w_014_018, w_005_038, w_005_046);
  and2 I014_020(w_014_020, w_009_202, w_009_027);
  nand2 I014_022(w_014_022, w_012_261, w_002_027);
  and2 I014_023(w_014_023, w_003_091, w_005_169);
  nand2 I014_024(w_014_024, w_013_044, w_005_115);
  or2  I014_025(w_014_025, w_009_020, w_013_215);
  and2 I014_027(w_014_027, w_003_019, w_012_016);
  or2  I014_028(w_014_028, w_004_132, w_006_000);
  or2  I014_033(w_014_033, w_005_200, w_003_042);
  nand2 I014_034(w_014_034, w_001_006, w_003_089);
  not1 I014_035(w_014_035, w_009_064);
  or2  I014_037(w_014_037, w_012_222, w_012_043);
  not1 I014_038(w_014_038, w_006_000);
  or2  I014_039(w_014_039, w_012_036, w_010_391);
  and2 I014_040(w_014_040, w_013_091, w_013_145);
  nand2 I014_043(w_014_043, w_005_065, w_006_000);
  and2 I014_044(w_014_044, w_002_015, w_006_000);
  or2  I014_045(w_014_045, w_011_317, w_012_249);
  or2  I014_046(w_014_046, w_009_140, w_001_006);
  nand2 I014_047(w_014_047, w_001_004, w_001_002);
  and2 I014_048(w_014_048, w_013_014, w_010_100);
  nand2 I014_049(w_014_049, w_001_001, w_001_002);
  nand2 I014_052(w_014_052, w_000_320, w_004_323);
  and2 I014_053(w_014_053, w_006_000, w_005_120);
  not1 I014_054(w_014_054, w_006_000);
  or2  I014_056(w_014_056, w_007_184, w_010_162);
  not1 I014_057(w_014_057, w_002_012);
  nand2 I014_058(w_014_058, w_010_152, w_001_001);
  not1 I014_059(w_014_059, w_008_125);
  not1 I014_060(w_014_060, w_008_180);
  nand2 I014_063(w_014_063, w_003_042, w_009_000);
  not1 I014_065(w_014_065, w_013_224);
  and2 I014_066(w_014_066, w_008_115, w_002_010);
  nand2 I014_067(w_014_067, w_002_020, w_002_012);
  or2  I014_068(w_014_068, w_006_000, w_007_298);
  or2  I014_069(w_014_069, w_002_020, w_013_054);
  nand2 I014_070(w_014_070, w_002_003, w_006_000);
  or2  I014_071(w_014_071, w_012_184, w_012_359);
  not1 I014_072(w_014_072, w_012_056);
  nand2 I014_073(w_014_073, w_001_004, w_004_137);
  or2  I014_074(w_014_074, w_004_373, w_004_137);
  nand2 I014_076(w_014_076, w_001_003, w_000_341);
  not1 I014_079(w_014_079, w_009_123);
  nand2 I014_080(w_014_080, w_012_260, w_001_003);
  or2  I014_081(w_014_081, w_003_089, w_010_449);
  and2 I014_082(w_014_082, w_012_339, w_007_027);
  and2 I014_083(w_014_083, w_006_000, w_012_097);
  and2 I014_084(w_014_084, w_002_016, w_007_006);
  not1 I014_085(w_014_085, w_005_052);
  and2 I014_086(w_014_086, w_013_159, w_012_357);
  and2 I014_087(w_014_087, w_013_217, w_003_056);
  nand2 I014_088(w_014_088, w_011_015, w_013_124);
  not1 I014_091(w_014_091, w_002_020);
  and2 I014_092(w_014_092, w_008_325, w_009_089);
  not1 I014_093(w_014_093, w_007_184);
  not1 I014_094(w_014_094, w_004_253);
  and2 I014_095(w_014_095, w_004_320, w_009_164);
  and2 I014_096(w_014_096, w_003_010, w_013_183);
  and2 I014_099(w_014_099, w_005_124, w_002_020);
  or2  I014_101(w_014_101, w_006_000, w_009_073);
  nand2 I014_102(w_014_102, w_004_327, w_007_273);
  or2  I014_103(w_014_103, w_004_457, w_003_046);
  or2  I014_104(w_014_104, w_004_036, w_005_034);
  and2 I014_105(w_014_105, w_000_326, w_009_084);
  not1 I014_106(w_014_106, w_006_000);
  and2 I014_108(w_014_108, w_005_192, w_008_245);
  and2 I014_109(w_014_109, w_013_019, w_009_152);
  and2 I014_110(w_014_110, w_011_196, w_007_391);
  nand2 I014_113(w_014_113, w_013_181, w_009_061);
  nand2 I014_114(w_014_114, w_001_002, w_012_050);
  not1 I014_115(w_014_115, w_008_309);
  or2  I014_116(w_014_116, w_003_097, w_013_080);
  or2  I014_118(w_014_118, w_004_004, w_005_235);
  and2 I014_119(w_014_119, w_004_061, w_003_075);
  or2  I014_121(w_014_121, w_001_002, w_013_142);
  and2 I014_122(w_014_122, w_000_368, w_005_192);
  or2  I014_123(w_014_123, w_011_000, w_006_000);
  not1 I014_125(w_014_125, w_012_116);
  or2  I014_128(w_014_128, w_013_176, w_006_000);
  and2 I014_129(w_014_129, w_011_163, w_001_002);
  or2  I014_131(w_014_131, w_000_411, w_001_005);
  nand2 I014_132(w_014_132, w_007_122, w_000_412);
  not1 I014_133(w_014_133, w_004_344);
  and2 I014_134(w_014_134, w_003_053, w_003_084);
  or2  I014_135(w_014_135, w_009_062, w_009_137);
  or2  I014_136(w_014_136, w_011_017, w_008_201);
  or2  I014_137(w_014_137, w_008_099, w_005_216);
  and2 I014_138(w_014_138, w_004_275, w_011_069);
  nand2 I014_140(w_014_140, w_009_107, w_010_417);
  nand2 I014_141(w_014_141, w_013_027, w_001_005);
  not1 I014_144(w_014_144, w_010_258);
  or2  I014_145(w_014_145, w_008_327, w_007_293);
  nand2 I014_146(w_014_146, w_006_000, w_012_298);
  nand2 I014_148(w_014_148, w_001_001, w_003_083);
  nand2 I014_150(w_014_150, w_012_040, w_013_168);
  not1 I014_151(w_014_151, w_006_000);
  or2  I014_152(w_014_152, w_011_051, w_002_020);
  nand2 I014_153(w_014_153, w_013_006, w_013_214);
  or2  I014_154(w_014_154, w_001_005, w_008_082);
  not1 I014_155(w_014_155, w_009_067);
  nand2 I014_156(w_014_156, w_003_083, w_010_294);
  and2 I014_157(w_014_157, w_006_000, w_003_093);
  or2  I014_159(w_014_159, w_010_349, w_012_090);
  or2  I014_161(w_014_161, w_003_019, w_007_154);
  and2 I014_163(w_014_163, w_001_002, w_008_153);
  and2 I014_164(w_014_164, w_010_445, w_008_104);
  nand2 I014_165(w_014_165, w_001_000, w_000_067);
  or2  I014_166(w_014_166, w_013_040, w_002_021);
  nand2 I014_167(w_014_167, w_013_187, w_013_081);
  and2 I014_169(w_014_169, w_001_004, w_006_000);
  not1 I014_170(w_014_170, w_000_028);
  and2 I014_173(w_014_173, w_007_121, w_009_020);
  or2  I014_174(w_014_174, w_006_000, w_004_089);
  nand2 I014_178(w_014_178, w_006_000, w_004_365);
  or2  I014_181(w_014_181, w_006_000, w_002_008);
  nand2 I014_182(w_014_182, w_013_038, w_009_089);
  or2  I014_183(w_014_183, w_012_042, w_009_059);
  nand2 I014_184(w_014_184, w_001_005, w_011_221);
  or2  I014_185(w_014_185, w_004_300, w_005_142);
  not1 I014_186(w_014_186, w_000_073);
  nand2 I014_188(w_014_188, w_009_194, w_006_000);
  not1 I014_191(w_014_191, w_005_023);
  not1 I014_193(w_014_193, w_011_134);
  nand2 I014_195(w_014_195, w_012_073, w_001_003);
  nand2 I014_196(w_014_196, w_007_316, w_004_211);
  and2 I014_197(w_014_197, w_004_001, w_010_054);
  and2 I014_198(w_014_198, w_002_005, w_013_226);
  and2 I014_202(w_014_202, w_011_095, w_004_395);
  not1 I014_203(w_014_203, w_007_072);
  not1 I014_204(w_014_204, w_001_004);
  not1 I014_205(w_014_205, w_001_002);
  or2  I014_206(w_014_206, w_008_325, w_008_228);
  nand2 I014_207(w_014_207, w_000_257, w_004_044);
  nand2 I014_208(w_014_208, w_011_334, w_001_000);
  and2 I014_209(w_014_209, w_010_333, w_009_137);
  or2  I014_210(w_014_210, w_010_038, w_008_146);
  or2  I014_211(w_014_211, w_007_030, w_013_122);
  nand2 I014_212(w_014_212, w_000_414, w_000_035);
  or2  I014_213(w_014_213, w_005_147, w_004_121);
  nand2 I014_215(w_014_215, w_006_000, w_004_083);
  nand2 I014_216(w_014_216, w_005_251, w_000_415);
  or2  I014_217(w_014_217, w_009_129, w_007_238);
  not1 I014_218(w_014_218, w_002_022);
  nand2 I014_219(w_014_219, w_001_001, w_011_234);
  or2  I014_220(w_014_220, w_013_208, w_007_325);
  not1 I014_221(w_014_221, w_001_000);
  or2  I014_222(w_014_222, w_007_383, w_011_113);
  and2 I014_225(w_014_225, w_007_261, w_005_011);
  and2 I014_226(w_014_226, w_006_000, w_005_008);
  not1 I014_227(w_014_227, w_005_216);
  nand2 I014_228(w_014_228, w_012_083, w_000_331);
  and2 I014_229(w_014_229, w_007_066, w_002_027);
  nand2 I014_231(w_014_231, w_011_035, w_012_024);
  or2  I014_233(w_014_233, w_009_233, w_001_000);
  not1 I014_234(w_014_234, w_002_017);
  or2  I014_235(w_014_235, w_002_016, w_001_005);
  nand2 I014_236(w_014_236, w_003_004, w_011_009);
  and2 I014_237(w_014_237, w_006_000, w_010_075);
  or2  I014_240(w_014_240, w_012_266, w_001_001);
  nand2 I014_241(w_014_241, w_010_018, w_008_000);
  not1 I014_243(w_014_243, w_007_386);
  or2  I014_245(w_014_245, w_005_013, w_002_026);
  nand2 I014_247(w_014_247, w_012_296, w_013_140);
  nand2 I014_248(w_014_248, w_011_084, w_008_087);
  and2 I014_249(w_014_249, w_004_340, w_003_099);
  and2 I014_252(w_014_252, w_003_008, w_010_048);
  not1 I014_254(w_014_254, w_010_451);
  not1 I014_256(w_014_256, w_000_240);
  not1 I014_259(w_014_259, w_011_088);
  or2  I014_260(w_014_260, w_010_429, w_011_093);
  not1 I014_262(w_014_262, w_010_034);
  not1 I014_264(w_014_264, w_008_010);
  not1 I014_265(w_014_265, w_000_104);
  not1 I015_000(w_015_000, w_007_063);
  nand2 I015_001(w_015_001, w_009_203, w_013_173);
  and2 I015_002(w_015_002, w_005_118, w_008_140);
  or2  I015_004(w_015_004, w_005_004, w_012_160);
  and2 I015_005(w_015_005, w_005_173, w_001_005);
  or2  I015_006(w_015_006, w_006_000, w_014_125);
  not1 I015_007(w_015_007, w_001_003);
  and2 I015_009(w_015_009, w_002_003, w_004_020);
  or2  I015_010(w_015_010, w_002_019, w_004_250);
  and2 I015_011(w_015_011, w_008_064, w_004_178);
  and2 I015_012(w_015_012, w_005_133, w_007_098);
  and2 I015_013(w_015_013, w_006_000, w_004_094);
  not1 I015_014(w_015_014, w_003_034);
  nand2 I015_015(w_015_015, w_004_137, w_000_296);
  and2 I015_017(w_015_017, w_002_026, w_008_119);
  and2 I015_018(w_015_018, w_004_021, w_002_023);
  not1 I015_020(w_015_020, w_000_225);
  and2 I015_021(w_015_021, w_000_416, w_012_225);
  nand2 I015_022(w_015_022, w_009_124, w_000_002);
  not1 I015_023(w_015_023, w_004_023);
  and2 I015_024(w_015_024, w_010_436, w_011_331);
  or2  I015_025(w_015_025, w_013_158, w_007_009);
  nand2 I015_026(w_015_026, w_008_243, w_013_011);
  or2  I015_027(w_015_027, w_014_006, w_008_103);
  not1 I015_028(w_015_028, w_005_026);
  or2  I015_029(w_015_029, w_006_000, w_009_151);
  not1 I015_031(w_015_031, w_005_201);
  and2 I015_033(w_015_033, w_011_054, w_013_032);
  nand2 I015_034(w_015_034, w_004_307, w_010_435);
  not1 I015_036(w_015_036, w_001_006);
  not1 I015_037(w_015_037, w_006_000);
  or2  I015_038(w_015_038, w_014_170, w_002_015);
  and2 I015_039(w_015_039, w_013_248, w_014_068);
  and2 I015_040(w_015_040, w_010_021, w_014_103);
  not1 I015_041(w_015_041, w_003_028);
  nand2 I015_042(w_015_042, w_013_205, w_002_021);
  or2  I015_043(w_015_043, w_009_199, w_006_000);
  or2  I015_044(w_015_044, w_012_057, w_014_216);
  not1 I015_045(w_015_045, w_008_083);
  not1 I015_046(w_015_046, w_006_000);
  and2 I015_047(w_015_047, w_006_000, w_000_261);
  not1 I015_048(w_015_048, w_004_395);
  not1 I015_049(w_015_049, w_004_234);
  not1 I015_050(w_015_050, w_003_074);
  nand2 I015_051(w_015_051, w_008_210, w_004_369);
  or2  I015_052(w_015_052, w_014_110, w_006_000);
  and2 I015_053(w_015_053, w_007_063, w_002_019);
  or2  I015_054(w_015_054, w_007_082, w_010_290);
  nand2 I015_055(w_015_055, w_013_132, w_013_075);
  not1 I015_058(w_015_058, w_012_091);
  nand2 I015_059(w_015_059, w_011_320, w_007_056);
  and2 I015_060(w_015_060, w_006_000, w_004_011);
  or2  I015_061(w_015_061, w_011_131, w_012_113);
  or2  I015_062(w_015_062, w_011_137, w_014_128);
  nand2 I015_063(w_015_063, w_009_052, w_014_169);
  not1 I015_064(w_015_064, w_007_391);
  and2 I015_065(w_015_065, w_011_335, w_008_047);
  nand2 I015_066(w_015_066, w_000_360, w_001_005);
  and2 I015_067(w_015_067, w_012_040, w_001_005);
  not1 I015_068(w_015_068, w_013_053);
  and2 I015_069(w_015_069, w_001_002, w_001_004);
  not1 I015_070(w_015_070, w_002_021);
  or2  I015_071(w_015_071, w_001_005, w_010_002);
  and2 I015_072(w_015_072, w_006_000, w_008_102);
  or2  I015_073(w_015_073, w_001_006, w_012_325);
  and2 I015_074(w_015_074, w_010_217, w_012_366);
  and2 I015_075(w_015_075, w_003_086, w_006_000);
  not1 I015_077(w_015_077, w_002_007);
  not1 I015_078(w_015_078, w_012_382);
  nand2 I015_080(w_015_080, w_009_025, w_009_002);
  not1 I015_081(w_015_081, w_001_006);
  not1 I015_082(w_015_082, w_003_086);
  and2 I015_083(w_015_083, w_014_243, w_006_000);
  not1 I015_085(w_015_085, w_007_124);
  not1 I015_086(w_015_086, w_007_264);
  not1 I015_088(w_015_088, w_011_088);
  and2 I015_089(w_015_089, w_004_359, w_004_246);
  and2 I015_090(w_015_090, w_004_302, w_011_182);
  nand2 I015_091(w_015_091, w_002_018, w_011_055);
  nand2 I015_092(w_015_092, w_001_006, w_013_013);
  and2 I015_093(w_015_093, w_005_024, w_004_020);
  and2 I015_095(w_015_095, w_009_078, w_014_220);
  or2  I015_096(w_015_096, w_010_014, w_004_419);
  or2  I015_097(w_015_097, w_001_005, w_005_142);
  nand2 I015_098(w_015_098, w_001_002, w_010_100);
  not1 I015_100(w_015_100, w_002_024);
  nand2 I015_102(w_015_102, w_000_239, w_005_064);
  or2  I015_105(w_015_105, w_004_015, w_012_159);
  not1 I015_106(w_015_106, w_012_272);
  not1 I015_108(w_015_108, w_014_146);
  or2  I015_111(w_015_111, w_013_084, w_010_103);
  or2  I015_112(w_015_112, w_000_093, w_000_276);
  nand2 I015_113(w_015_113, w_012_049, w_013_052);
  nand2 I015_114(w_015_114, w_005_214, w_001_002);
  nand2 I015_115(w_015_115, w_000_410, w_004_189);
  not1 I015_116(w_015_116, w_005_038);
  and2 I015_117(w_015_117, w_001_006, w_006_000);
  or2  I015_120(w_015_120, w_006_000, w_001_004);
  or2  I015_121(w_015_121, w_006_000, w_005_043);
  not1 I015_122(w_015_122, w_005_052);
  nand2 I015_124(w_015_124, w_001_006, w_010_441);
  or2  I015_125(w_015_125, w_012_366, w_010_196);
  and2 I015_126(w_015_126, w_004_416, w_010_062);
  not1 I015_127(w_015_127, w_011_111);
  nand2 I015_128(w_015_128, w_009_223, w_003_000);
  nand2 I015_129(w_015_129, w_000_213, w_002_003);
  nand2 I015_131(w_015_131, w_000_107, w_006_000);
  or2  I015_132(w_015_132, w_008_139, w_000_412);
  and2 I015_134(w_015_134, w_013_012, w_000_417);
  and2 I016_001(w_016_001, w_011_153, w_006_000);
  nand2 I016_002(w_016_002, w_009_113, w_004_362);
  nand2 I016_003(w_016_003, w_014_072, w_008_072);
  nand2 I016_005(w_016_005, w_009_000, w_004_011);
  and2 I016_007(w_016_007, w_006_000, w_010_204);
  nand2 I016_008(w_016_008, w_001_002, w_014_221);
  and2 I016_009(w_016_009, w_005_039, w_004_113);
  and2 I016_011(w_016_011, w_010_372, w_010_318);
  and2 I016_012(w_016_012, w_006_000, w_003_048);
  nand2 I016_014(w_016_014, w_010_223, w_012_001);
  and2 I016_015(w_016_015, w_004_314, w_000_217);
  nand2 I016_016(w_016_016, w_015_054, w_000_418);
  or2  I016_017(w_016_017, w_012_277, w_006_000);
  and2 I016_018(w_016_018, w_010_441, w_013_109);
  or2  I016_019(w_016_019, w_012_010, w_011_028);
  nand2 I016_020(w_016_020, w_002_010, w_006_000);
  nand2 I016_021(w_016_021, w_003_055, w_009_231);
  and2 I016_022(w_016_022, w_004_178, w_010_035);
  or2  I016_023(w_016_023, w_000_217, w_011_254);
  and2 I016_024(w_016_024, w_011_133, w_005_112);
  or2  I016_026(w_016_026, w_006_000, w_015_021);
  nand2 I016_027(w_016_027, w_010_404, w_006_000);
  nand2 I016_028(w_016_028, w_003_022, w_005_208);
  and2 I016_029(w_016_029, w_015_081, w_013_229);
  nand2 I016_030(w_016_030, w_005_177, w_003_000);
  or2  I016_031(w_016_031, w_001_005, w_002_012);
  not1 I016_032(w_016_032, w_015_002);
  not1 I016_033(w_016_033, w_015_011);
  or2  I016_034(w_016_034, w_009_051, w_015_045);
  not1 I016_035(w_016_035, w_002_005);
  nand2 I016_037(w_016_037, w_013_200, w_004_350);
  and2 I016_038(w_016_038, w_015_083, w_005_206);
  or2  I016_044(w_016_044, w_001_000, w_005_012);
  nand2 I016_045(w_016_045, w_011_128, w_009_022);
  or2  I016_046(w_016_046, w_010_120, w_008_085);
  and2 I016_048(w_016_048, w_000_247, w_008_142);
  not1 I016_049(w_016_049, w_005_118);
  nand2 I016_051(w_016_051, w_003_063, w_004_159);
  not1 I016_052(w_016_052, w_015_074);
  nand2 I016_053(w_016_053, w_008_243, w_006_000);
  not1 I016_056(w_016_056, w_014_235);
  and2 I016_058(w_016_058, w_004_224, w_009_009);
  not1 I016_059(w_016_059, w_008_082);
  and2 I016_061(w_016_061, w_013_169, w_001_003);
  not1 I016_062(w_016_062, w_007_309);
  and2 I016_065(w_016_065, w_000_179, w_008_126);
  and2 I016_067(w_016_067, w_009_147, w_004_454);
  or2  I016_068(w_016_068, w_005_028, w_015_064);
  and2 I016_070(w_016_070, w_001_001, w_011_125);
  not1 I016_071(w_016_071, w_015_080);
  not1 I016_073(w_016_073, w_007_347);
  nand2 I016_074(w_016_074, w_001_002, w_013_113);
  or2  I016_076(w_016_076, w_002_008, w_005_126);
  not1 I016_077(w_016_077, w_007_276);
  nand2 I016_078(w_016_078, w_007_082, w_008_089);
  not1 I016_079(w_016_079, w_008_283);
  or2  I016_080(w_016_080, w_005_133, w_009_204);
  nand2 I016_082(w_016_082, w_002_025, w_013_088);
  and2 I016_084(w_016_084, w_004_322, w_008_045);
  or2  I016_085(w_016_085, w_000_420, w_011_332);
  and2 I016_086(w_016_086, w_013_189, w_006_000);
  or2  I016_087(w_016_087, w_007_032, w_001_001);
  and2 I016_091(w_016_091, w_003_010, w_008_068);
  or2  I016_093(w_016_093, w_011_091, w_002_020);
  and2 I016_094(w_016_094, w_006_000, w_012_127);
  not1 I016_095(w_016_095, w_005_080);
  not1 I016_097(w_016_097, w_011_289);
  not1 I016_099(w_016_099, w_013_197);
  nand2 I016_101(w_016_101, w_015_012, w_003_009);
  not1 I016_106(w_016_106, w_009_137);
  nand2 I016_107(w_016_107, w_002_016, w_011_143);
  or2  I016_110(w_016_110, w_004_157, w_006_000);
  nand2 I016_111(w_016_111, w_005_065, w_006_000);
  or2  I016_113(w_016_113, w_002_021, w_013_094);
  and2 I016_117(w_016_117, w_000_317, w_014_080);
  not1 I016_118(w_016_118, w_007_380);
  not1 I016_119(w_016_119, w_007_019);
  and2 I016_122(w_016_122, w_005_217, w_008_039);
  nand2 I016_124(w_016_124, w_010_317, w_015_015);
  nand2 I016_125(w_016_125, w_005_000, w_015_045);
  not1 I016_130(w_016_130, w_014_210);
  and2 I016_133(w_016_133, w_008_001, w_002_001);
  or2  I016_136(w_016_136, w_010_268, w_011_164);
  or2  I016_139(w_016_139, w_015_048, w_012_042);
  and2 I016_140(w_016_140, w_004_389, w_002_025);
  and2 I016_141(w_016_141, w_004_043, w_006_000);
  not1 I016_144(w_016_144, w_004_407);
  not1 I016_145(w_016_145, w_006_000);
  and2 I016_147(w_016_147, w_006_000, w_012_039);
  not1 I016_149(w_016_149, w_006_000);
  or2  I016_151(w_016_151, w_000_261, w_003_079);
  not1 I016_152(w_016_152, w_010_024);
  and2 I016_153(w_016_153, w_013_112, w_014_025);
  or2  I016_157(w_016_157, w_009_115, w_006_000);
  and2 I016_164(w_016_164, w_013_065, w_001_003);
  nand2 I016_165(w_016_165, w_002_001, w_006_000);
  not1 I016_169(w_016_169, w_004_225);
  and2 I016_173(w_016_173, w_010_362, w_005_123);
  not1 I016_175(w_016_175, w_013_134);
  or2  I016_176(w_016_176, w_001_004, w_010_328);
  not1 I016_177(w_016_177, w_003_070);
  or2  I016_178(w_016_178, w_013_243, w_007_017);
  or2  I016_182(w_016_182, w_011_077, w_002_013);
  and2 I016_183(w_016_183, w_012_261, w_010_030);
  nand2 I016_185(w_016_185, w_011_132, w_005_065);
  and2 I016_187(w_016_187, w_006_000, w_007_068);
  or2  I016_189(w_016_189, w_006_000, w_010_180);
  nand2 I016_191(w_016_191, w_003_041, w_014_069);
  or2  I016_192(w_016_192, w_005_001, w_005_229);
  nand2 I016_194(w_016_194, w_001_004, w_004_023);
  or2  I016_197(w_016_197, w_001_002, w_002_021);
  not1 I016_200(w_016_200, w_005_149);
  and2 I016_209(w_016_209, w_013_062, w_008_156);
  not1 I016_210(w_016_210, w_000_422);
  nand2 I016_212(w_016_212, w_014_159, w_013_210);
  nand2 I016_213(w_016_213, w_002_010, w_010_412);
  and2 I016_214(w_016_214, w_013_147, w_000_078);
  not1 I016_216(w_016_216, w_005_023);
  not1 I016_222(w_016_222, w_011_204);
  nand2 I016_223(w_016_223, w_010_343, w_004_173);
  and2 I016_225(w_016_225, w_011_177, w_008_150);
  or2  I016_228(w_016_228, w_008_275, w_002_010);
  not1 I016_230(w_016_230, w_008_234);
  not1 I016_232(w_016_232, w_011_023);
  not1 I016_233(w_016_233, w_006_000);
  and2 I016_234(w_016_234, w_006_000, w_010_044);
  not1 I016_239(w_016_239, w_012_028);
  nand2 I016_241(w_016_241, w_007_321, w_011_090);
  nand2 I016_244(w_016_244, w_012_322, w_003_077);
  or2  I016_245(w_016_245, w_004_178, w_007_308);
  nand2 I016_247(w_016_247, w_001_003, w_007_340);
  nand2 I016_248(w_016_248, w_002_011, w_006_000);
  nand2 I016_249(w_016_249, w_002_020, w_015_048);
  nand2 I016_250(w_016_250, w_011_142, w_014_056);
  and2 I016_253(w_016_253, w_009_021, w_002_000);
  or2  I016_254(w_016_254, w_002_002, w_004_152);
  and2 I016_255(w_016_255, w_000_138, w_000_071);
  not1 I016_256(w_016_256, w_012_147);
  nand2 I016_257(w_016_257, w_010_055, w_010_384);
  and2 I016_258(w_016_258, w_015_054, w_015_083);
  and2 I016_260(w_016_260, w_003_050, w_005_068);
  and2 I016_262(w_016_262, w_001_006, w_002_009);
  and2 I016_263(w_016_263, w_006_000, w_007_376);
  and2 I016_264(w_016_264, w_003_019, w_007_019);
  not1 I016_265(w_016_265, w_015_108);
  or2  I016_268(w_016_268, w_005_235, w_013_046);
  not1 I016_274(w_016_274, w_005_027);
  and2 I016_278(w_016_278, w_012_191, w_008_191);
  not1 I016_279(w_016_279, w_014_207);
  nand2 I016_280(w_016_280, w_006_000, w_008_038);
  and2 I016_281(w_016_281, w_014_264, w_000_257);
  and2 I016_285(w_016_285, w_004_166, w_009_012);
  and2 I016_286(w_016_286, w_007_071, w_004_285);
  and2 I016_287(w_016_287, w_012_170, w_000_398);
  and2 I016_291(w_016_291, w_013_199, w_000_125);
  not1 I016_292(w_016_292, w_009_013);
  not1 I016_294(w_016_294, w_014_131);
  nand2 I016_295(w_016_295, w_000_365, w_005_013);
  and2 I016_297(w_016_297, w_007_064, w_013_027);
  not1 I016_300(w_016_300, w_004_078);
  nand2 I016_301(w_016_301, w_000_345, w_014_011);
  or2  I016_303(w_016_303, w_010_036, w_013_162);
  or2  I016_304(w_016_304, w_010_189, w_001_004);
  nand2 I016_310(w_016_310, w_004_054, w_004_366);
  and2 I016_311(w_016_311, w_010_201, w_007_108);
  not1 I016_315(w_016_315, w_013_208);
  not1 I016_316(w_016_316, w_012_146);
  not1 I016_319(w_016_319, w_012_109);
  nand2 I016_322(w_016_322, w_005_133, w_004_070);
  or2  I016_324(w_016_324, w_015_022, w_015_127);
  not1 I016_328(w_016_328, w_007_388);
  nand2 I016_330(w_016_330, w_002_019, w_009_043);
  or2  I016_335(w_016_335, w_004_457, w_005_111);
  and2 I016_336(w_016_336, w_014_202, w_008_092);
  or2  I016_337(w_016_337, w_001_002, w_006_000);
  and2 I016_339(w_016_339, w_011_004, w_008_117);
  not1 I016_345(w_016_345, w_003_008);
  not1 I016_347(w_016_347, w_010_214);
  and2 I016_349(w_016_349, w_005_184, w_008_152);
  or2  I016_350(w_016_350, w_006_000, w_015_011);
  or2  I016_354(w_016_354, w_008_291, w_011_123);
  and2 I016_355(w_016_355, w_012_097, w_012_012);
  and2 I016_356(w_016_356, w_002_016, w_004_118);
  or2  I016_357(w_016_357, w_011_026, w_012_350);
  nand2 I016_362(w_016_362, w_009_074, w_003_019);
  nand2 I016_364(w_016_364, w_003_062, w_011_337);
  nand2 I016_367(w_016_367, w_005_162, w_014_011);
  nand2 I016_369(w_016_369, w_012_019, w_015_023);
  not1 I016_371(w_016_371, w_006_000);
  nand2 I016_372(w_016_372, w_014_054, w_005_010);
  nand2 I016_374(w_016_374, w_006_000, w_003_086);
  nand2 I016_375(w_016_375, w_014_084, w_005_088);
  or2  I016_378(w_016_378, w_002_005, w_008_008);
  or2  I016_380(w_016_380, w_012_318, w_000_425);
  or2  I016_381(w_016_381, w_007_206, w_004_017);
  not1 I016_382(w_016_382, w_002_003);
  and2 I016_384(w_016_384, w_005_171, w_001_001);
  and2 I016_385(w_016_385, w_009_148, w_000_135);
  nand2 I016_391(w_016_391, w_007_245, w_003_059);
  not1 I016_394(w_016_394, w_010_240);
  or2  I016_395(w_016_395, w_014_136, w_010_265);
  not1 I016_398(w_016_398, w_013_006);
  not1 I016_399(w_016_399, w_005_008);
  not1 I017_000(w_017_000, w_014_053);
  not1 I017_001(w_017_001, w_013_017);
  or2  I017_003(w_017_003, w_013_044, w_009_121);
  nand2 I017_004(w_017_004, w_015_124, w_001_000);
  not1 I017_005(w_017_005, w_005_201);
  not1 I017_006(w_017_006, w_015_067);
  and2 I017_007(w_017_007, w_014_033, w_014_056);
  not1 I017_008(w_017_008, w_006_000);
  or2  I017_009(w_017_009, w_002_022, w_015_059);
  and2 I017_010(w_017_010, w_001_005, w_004_460);
  and2 I017_011(w_017_011, w_000_219, w_008_075);
  nand2 I017_012(w_017_012, w_004_008, w_015_038);
  not1 I017_014(w_017_014, w_009_161);
  nand2 I017_015(w_017_015, w_015_078, w_012_186);
  nand2 I017_016(w_017_016, w_006_000, w_003_044);
  and2 I017_017(w_017_017, w_012_045, w_007_125);
  and2 I017_018(w_017_018, w_015_072, w_001_001);
  nand2 I017_019(w_017_019, w_013_054, w_010_211);
  or2  I017_020(w_017_020, w_005_077, w_015_097);
  and2 I017_021(w_017_021, w_004_406, w_005_119);
  and2 I017_022(w_017_022, w_010_364, w_009_088);
  and2 I017_023(w_017_023, w_012_253, w_015_009);
  not1 I017_024(w_017_024, w_000_174);
  not1 I017_025(w_017_025, w_010_137);
  not1 I017_026(w_017_026, w_006_000);
  not1 I017_027(w_017_027, w_014_203);
  and2 I017_028(w_017_028, w_002_000, w_001_001);
  not1 I017_029(w_017_029, w_005_148);
  not1 I017_030(w_017_030, w_010_218);
  or2  I017_033(w_017_033, w_009_221, w_010_037);
  or2  I017_034(w_017_034, w_015_004, w_016_260);
  and2 I017_035(w_017_035, w_001_001, w_009_189);
  not1 I017_036(w_017_036, w_014_074);
  or2  I017_037(w_017_037, w_015_068, w_008_079);
  not1 I017_038(w_017_038, w_001_006);
  or2  I017_039(w_017_039, w_007_001, w_005_088);
  not1 I017_040(w_017_040, w_015_029);
  not1 I017_041(w_017_041, w_008_250);
  and2 I017_042(w_017_042, w_000_363, w_009_104);
  not1 I017_043(w_017_043, w_000_244);
  not1 I017_044(w_017_044, w_009_104);
  and2 I017_045(w_017_045, w_014_198, w_001_003);
  nand2 I017_046(w_017_046, w_011_034, w_012_380);
  not1 I017_047(w_017_047, w_010_101);
  and2 I017_048(w_017_048, w_007_200, w_002_011);
  not1 I017_049(w_017_049, w_012_275);
  nand2 I017_050(w_017_050, w_004_324, w_016_145);
  or2  I017_051(w_017_051, w_014_105, w_011_058);
  nand2 I017_052(w_017_052, w_008_020, w_005_021);
  or2  I017_053(w_017_053, w_007_160, w_016_301);
  not1 I017_054(w_017_054, w_009_165);
  not1 I017_055(w_017_055, w_008_109);
  nand2 I017_056(w_017_056, w_005_097, w_016_015);
  and2 I017_058(w_017_058, w_010_077, w_005_153);
  and2 I017_059(w_017_059, w_005_118, w_010_219);
  or2  I017_060(w_017_060, w_008_231, w_007_025);
  or2  I017_061(w_017_061, w_008_185, w_005_009);
  and2 I017_063(w_017_063, w_009_115, w_003_001);
  or2  I017_064(w_017_064, w_005_000, w_013_113);
  nand2 I017_065(w_017_065, w_001_002, w_002_017);
  or2  I017_066(w_017_066, w_010_389, w_012_056);
  nand2 I017_067(w_017_067, w_014_229, w_014_265);
  nand2 I017_070(w_017_070, w_008_118, w_004_309);
  nand2 I017_071(w_017_071, w_003_011, w_005_130);
  and2 I017_072(w_017_072, w_013_246, w_015_074);
  or2  I017_073(w_017_073, w_006_000, w_007_337);
  or2  I017_074(w_017_074, w_006_000, w_000_397);
  or2  I017_075(w_017_075, w_001_001, w_013_055);
  and2 I017_076(w_017_076, w_012_262, w_014_228);
  nand2 I017_077(w_017_077, w_003_024, w_003_080);
  not1 I017_078(w_017_078, w_000_304);
  or2  I017_080(w_017_080, w_001_004, w_013_061);
  and2 I017_081(w_017_081, w_013_189, w_010_193);
  not1 I017_083(w_017_083, w_009_120);
  or2  I017_084(w_017_084, w_003_042, w_007_106);
  nand2 I017_085(w_017_085, w_015_002, w_003_033);
  and2 I017_086(w_017_086, w_006_000, w_007_228);
  and2 I017_087(w_017_087, w_006_000, w_003_040);
  not1 I017_088(w_017_088, w_004_047);
  or2  I017_091(w_017_091, w_014_237, w_006_000);
  nand2 I017_092(w_017_092, w_000_168, w_000_426);
  not1 I017_093(w_017_093, w_015_039);
  or2  I017_094(w_017_094, w_009_033, w_005_192);
  and2 I017_098(w_017_098, w_006_000, w_014_071);
  or2  I017_099(w_017_099, w_006_000, w_007_196);
  or2  I017_100(w_017_100, w_005_118, w_002_015);
  not1 I017_101(w_017_101, w_015_128);
  not1 I017_103(w_017_103, w_014_034);
  or2  I017_104(w_017_104, w_013_265, w_010_072);
  nand2 I017_108(w_017_108, w_004_430, w_014_161);
  or2  I017_109(w_017_109, w_007_221, w_013_213);
  and2 I017_111(w_017_111, w_004_357, w_004_128);
  and2 I017_113(w_017_113, w_003_063, w_013_102);
  not1 I017_114(w_017_114, w_011_058);
  and2 I017_115(w_017_115, w_008_062, w_008_161);
  nand2 I017_116(w_017_116, w_004_374, w_006_000);
  and2 I017_117(w_017_117, w_012_282, w_011_097);
  nand2 I017_118(w_017_118, w_015_068, w_012_293);
  nand2 I017_122(w_017_122, w_008_054, w_012_313);
  and2 I017_123(w_017_123, w_007_188, w_010_311);
  and2 I017_124(w_017_124, w_005_192, w_005_006);
  and2 I017_126(w_017_126, w_004_066, w_011_297);
  or2  I017_128(w_017_128, w_013_008, w_012_225);
  or2  I017_130(w_017_130, w_015_077, w_004_115);
  and2 I017_133(w_017_133, w_001_001, w_001_003);
  not1 I017_135(w_017_135, w_005_194);
  nand2 I017_136(w_017_136, w_005_212, w_003_083);
  or2  I017_138(w_017_138, w_011_127, w_016_056);
  and2 I017_139(w_017_139, w_004_426, w_010_264);
  or2  I017_141(w_017_141, w_013_199, w_013_039);
  or2  I017_143(w_017_143, w_006_000, w_015_045);
  and2 I017_144(w_017_144, w_015_068, w_000_196);
  not1 I017_146(w_017_146, w_012_030);
  or2  I017_148(w_017_148, w_011_153, w_002_010);
  not1 I017_150(w_017_150, w_008_124);
  and2 I017_154(w_017_154, w_001_004, w_009_186);
  nand2 I017_155(w_017_155, w_004_430, w_004_241);
  nand2 I017_156(w_017_156, w_008_310, w_005_049);
  and2 I017_157(w_017_157, w_013_009, w_011_318);
  nand2 I017_159(w_017_159, w_012_131, w_003_092);
  and2 I017_162(w_017_162, w_005_049, w_007_299);
  and2 I017_163(w_017_163, w_000_427, w_014_024);
  and2 I017_166(w_017_166, w_003_094, w_002_006);
  and2 I017_167(w_017_167, w_012_030, w_003_026);
  or2  I017_168(w_017_168, w_003_088, w_003_044);
  nand2 I017_171(w_017_171, w_008_337, w_010_188);
  not1 I017_172(w_017_172, w_005_136);
  nand2 I017_173(w_017_173, w_015_134, w_012_084);
  nand2 I017_176(w_017_176, w_000_389, w_001_001);
  or2  I017_177(w_017_177, w_010_267, w_001_006);
  and2 I017_178(w_017_178, w_002_005, w_009_204);
  not1 I017_179(w_017_179, w_010_224);
  and2 I017_180(w_017_180, w_013_161, w_009_104);
  nand2 I017_181(w_017_181, w_012_030, w_009_072);
  nand2 I017_182(w_017_182, w_016_264, w_004_199);
  nand2 I017_184(w_017_184, w_014_045, w_009_075);
  and2 I017_185(w_017_185, w_012_295, w_014_099);
  or2  I017_186(w_017_186, w_007_176, w_008_000);
  or2  I017_187(w_017_187, w_001_005, w_012_186);
  nand2 I017_188(w_017_188, w_005_006, w_016_304);
  nand2 I017_190(w_017_190, w_001_004, w_001_006);
  nand2 I017_191(w_017_191, w_006_000, w_003_050);
  nand2 I018_000(w_018_000, w_001_000, w_015_073);
  or2  I018_001(w_018_001, w_014_113, w_008_040);
  and2 I018_002(w_018_002, w_015_089, w_014_025);
  or2  I018_003(w_018_003, w_010_381, w_016_152);
  not1 I018_005(w_018_005, w_002_016);
  and2 I018_006(w_018_006, w_002_000, w_014_191);
  not1 I018_008(w_018_008, w_000_143);
  or2  I018_010(w_018_010, w_017_014, w_017_020);
  and2 I018_012(w_018_012, w_008_110, w_010_398);
  and2 I018_014(w_018_014, w_002_003, w_002_023);
  or2  I018_015(w_018_015, w_001_004, w_003_050);
  nand2 I018_016(w_018_016, w_012_039, w_013_047);
  nand2 I018_017(w_018_017, w_000_220, w_008_345);
  not1 I018_018(w_018_018, w_016_012);
  nand2 I018_019(w_018_019, w_008_064, w_000_397);
  or2  I018_020(w_018_020, w_009_008, w_017_155);
  and2 I018_022(w_018_022, w_001_005, w_008_184);
  nand2 I018_023(w_018_023, w_001_000, w_000_429);
  not1 I018_026(w_018_026, w_010_134);
  or2  I018_027(w_018_027, w_015_098, w_003_033);
  or2  I018_030(w_018_030, w_011_117, w_002_027);
  nand2 I018_031(w_018_031, w_017_033, w_002_018);
  not1 I018_032(w_018_032, w_015_031);
  and2 I018_034(w_018_034, w_016_084, w_006_000);
  or2  I018_035(w_018_035, w_001_001, w_014_259);
  not1 I018_037(w_018_037, w_008_264);
  not1 I018_039(w_018_039, w_006_000);
  or2  I018_040(w_018_040, w_007_372, w_001_004);
  not1 I018_045(w_018_045, w_010_123);
  nand2 I018_047(w_018_047, w_000_277, w_009_192);
  and2 I018_048(w_018_048, w_017_043, w_016_026);
  not1 I018_050(w_018_050, w_013_182);
  nand2 I018_051(w_018_051, w_014_023, w_016_008);
  or2  I018_053(w_018_053, w_010_065, w_008_261);
  not1 I018_054(w_018_054, w_015_033);
  nand2 I018_057(w_018_057, w_016_356, w_003_026);
  and2 I018_059(w_018_059, w_010_035, w_007_134);
  not1 I018_060(w_018_060, w_016_395);
  and2 I018_061(w_018_061, w_011_200, w_015_028);
  nand2 I018_063(w_018_063, w_012_015, w_002_014);
  not1 I018_064(w_018_064, w_005_052);
  and2 I018_067(w_018_067, w_003_097, w_016_027);
  nand2 I018_068(w_018_068, w_007_078, w_007_360);
  or2  I018_070(w_018_070, w_009_021, w_009_003);
  not1 I018_071(w_018_071, w_013_024);
  or2  I018_072(w_018_072, w_013_126, w_012_103);
  not1 I018_074(w_018_074, w_001_001);
  and2 I018_075(w_018_075, w_014_123, w_011_041);
  and2 I018_076(w_018_076, w_005_172, w_002_025);
  not1 I018_078(w_018_078, w_002_010);
  not1 I018_080(w_018_080, w_004_267);
  not1 I018_081(w_018_081, w_001_003);
  and2 I018_083(w_018_083, w_000_405, w_000_406);
  or2  I018_084(w_018_084, w_001_004, w_000_216);
  or2  I018_086(w_018_086, w_013_028, w_015_014);
  nand2 I018_089(w_018_089, w_016_330, w_005_149);
  or2  I018_091(w_018_091, w_011_253, w_011_083);
  and2 I018_094(w_018_094, w_007_219, w_010_410);
  and2 I018_095(w_018_095, w_017_036, w_016_009);
  nand2 I018_096(w_018_096, w_011_081, w_017_118);
  or2  I018_097(w_018_097, w_017_018, w_008_206);
  and2 I018_098(w_018_098, w_007_214, w_004_014);
  and2 I018_100(w_018_100, w_014_017, w_015_102);
  or2  I018_102(w_018_102, w_013_090, w_015_052);
  or2  I018_103(w_018_103, w_011_110, w_007_053);
  nand2 I018_104(w_018_104, w_000_235, w_004_460);
  and2 I018_105(w_018_105, w_010_306, w_007_389);
  not1 I018_106(w_018_106, w_016_337);
  or2  I018_107(w_018_107, w_011_064, w_004_159);
  and2 I018_108(w_018_108, w_012_364, w_011_001);
  nand2 I018_110(w_018_110, w_002_015, w_003_038);
  not1 I018_111(w_018_111, w_005_157);
  not1 I018_112(w_018_112, w_015_055);
  not1 I018_114(w_018_114, w_006_000);
  not1 I018_118(w_018_118, w_006_000);
  not1 I018_119(w_018_119, w_010_384);
  or2  I018_123(w_018_123, w_013_084, w_006_000);
  not1 I018_124(w_018_124, w_013_103);
  or2  I018_125(w_018_125, w_006_000, w_011_066);
  and2 I018_126(w_018_126, w_001_000, w_003_066);
  or2  I018_127(w_018_127, w_004_238, w_003_057);
  nand2 I018_130(w_018_130, w_005_066, w_010_020);
  or2  I018_131(w_018_131, w_003_020, w_012_099);
  not1 I018_132(w_018_132, w_006_000);
  not1 I018_133(w_018_133, w_007_007);
  or2  I018_134(w_018_134, w_003_000, w_000_074);
  not1 I018_135(w_018_135, w_003_019);
  or2  I018_136(w_018_136, w_011_280, w_017_139);
  or2  I018_137(w_018_137, w_002_022, w_000_181);
  and2 I018_139(w_018_139, w_004_312, w_001_003);
  and2 I018_141(w_018_141, w_017_167, w_009_126);
  nand2 I018_142(w_018_142, w_011_226, w_000_336);
  nand2 I018_143(w_018_143, w_011_116, w_012_358);
  not1 I018_144(w_018_144, w_013_105);
  not1 I018_145(w_018_145, w_006_000);
  and2 I018_146(w_018_146, w_006_000, w_002_010);
  and2 I018_150(w_018_150, w_003_091, w_017_155);
  or2  I018_151(w_018_151, w_012_260, w_015_112);
  and2 I018_153(w_018_153, w_012_219, w_005_073);
  and2 I018_155(w_018_155, w_004_273, w_001_003);
  nand2 I018_156(w_018_156, w_005_151, w_006_000);
  and2 I018_157(w_018_157, w_017_038, w_010_235);
  not1 I018_158(w_018_158, w_008_140);
  nand2 I018_160(w_018_160, w_006_000, w_011_150);
  or2  I018_161(w_018_161, w_006_000, w_013_184);
  or2  I018_162(w_018_162, w_012_291, w_012_088);
  and2 I018_163(w_018_163, w_017_070, w_014_122);
  or2  I018_164(w_018_164, w_006_000, w_005_052);
  and2 I018_165(w_018_165, w_002_009, w_002_005);
  and2 I018_167(w_018_167, w_017_128, w_004_107);
  and2 I018_168(w_018_168, w_013_141, w_006_000);
  or2  I018_169(w_018_169, w_010_241, w_002_004);
  or2  I018_171(w_018_171, w_009_160, w_010_317);
  nand2 I018_173(w_018_173, w_013_018, w_017_130);
  and2 I018_175(w_018_175, w_006_000, w_001_005);
  nand2 I018_181(w_018_181, w_012_180, w_013_225);
  and2 I018_182(w_018_182, w_007_234, w_006_000);
  and2 I018_183(w_018_183, w_002_005, w_005_164);
  nand2 I018_186(w_018_186, w_003_033, w_015_068);
  or2  I018_187(w_018_187, w_008_177, w_007_065);
  and2 I018_196(w_018_196, w_007_368, w_005_242);
  nand2 I018_197(w_018_197, w_003_015, w_003_040);
  or2  I018_199(w_018_199, w_014_086, w_001_000);
  or2  I018_200(w_018_200, w_004_163, w_008_106);
  not1 I018_203(w_018_203, w_015_000);
  and2 I018_206(w_018_206, w_003_096, w_007_222);
  and2 I018_211(w_018_211, w_002_015, w_003_074);
  or2  I018_212(w_018_212, w_010_226, w_001_000);
  or2  I018_213(w_018_213, w_006_000, w_013_149);
  and2 I018_215(w_018_215, w_000_172, w_006_000);
  or2  I018_218(w_018_218, w_013_186, w_001_003);
  and2 I018_229(w_018_229, w_010_012, w_002_002);
  and2 I018_234(w_018_234, w_004_142, w_012_097);
  nand2 I018_235(w_018_235, w_015_006, w_014_099);
  nand2 I018_236(w_018_236, w_016_068, w_007_090);
  nand2 I018_237(w_018_237, w_017_094, w_017_011);
  and2 I018_239(w_018_239, w_009_183, w_017_184);
  not1 I018_243(w_018_243, w_016_071);
  and2 I018_246(w_018_246, w_010_286, w_017_045);
  and2 I018_248(w_018_248, w_014_213, w_006_000);
  and2 I018_249(w_018_249, w_006_000, w_015_025);
  not1 I018_250(w_018_250, w_013_096);
  nand2 I018_256(w_018_256, w_016_065, w_016_144);
  not1 I018_257(w_018_257, w_005_236);
  or2  I018_259(w_018_259, w_009_196, w_008_068);
  not1 I018_263(w_018_263, w_009_125);
  or2  I018_270(w_018_270, w_016_044, w_009_104);
  nand2 I018_278(w_018_278, w_007_247, w_015_106);
  or2  I018_279(w_018_279, w_010_261, w_017_017);
  not1 I018_282(w_018_282, w_005_169);
  not1 I018_283(w_018_283, w_004_312);
  and2 I018_285(w_018_285, w_002_018, w_014_060);
  or2  I018_287(w_018_287, w_008_048, w_009_190);
  and2 I018_288(w_018_288, w_011_096, w_010_354);
  or2  I018_291(w_018_291, w_005_139, w_009_001);
  and2 I018_292(w_018_292, w_007_288, w_011_179);
  nand2 I018_293(w_018_293, w_005_152, w_010_362);
  or2  I018_295(w_018_295, w_000_352, w_012_028);
  not1 I018_297(w_018_297, w_013_245);
  nand2 I018_300(w_018_300, w_009_123, w_015_132);
  or2  I018_301(w_018_301, w_007_265, w_010_448);
  or2  I018_302(w_018_302, w_004_328, w_003_035);
  not1 I018_306(w_018_306, w_012_241);
  not1 I018_311(w_018_311, w_009_156);
  not1 I018_312(w_018_312, w_009_099);
  nand2 I018_313(w_018_313, w_012_176, w_002_020);
  or2  I018_314(w_018_314, w_011_150, w_017_016);
  and2 I018_320(w_018_320, w_002_016, w_011_181);
  or2  I018_321(w_018_321, w_006_000, w_010_159);
  not1 I018_322(w_018_322, w_001_004);
  nand2 I019_000(w_019_000, w_006_000, w_013_025);
  and2 I019_001(w_019_001, w_001_002, w_000_339);
  nand2 I019_002(w_019_002, w_005_077, w_016_212);
  not1 I019_003(w_019_003, w_013_228);
  not1 I019_004(w_019_004, w_007_126);
  and2 I019_005(w_019_005, w_015_075, w_004_376);
  not1 I019_006(w_019_006, w_000_379);
  or2  I019_007(w_019_007, w_010_255, w_004_109);
  not1 I019_008(w_019_008, w_006_000);
  not1 I019_009(w_019_009, w_014_227);
  or2  I019_010(w_019_010, w_008_223, w_003_060);
  nand2 I019_011(w_019_011, w_006_000, w_004_340);
  not1 I019_012(w_019_012, w_004_188);
  nand2 I019_013(w_019_013, w_004_446, w_002_016);
  not1 I019_014(w_019_014, w_003_077);
  and2 I019_015(w_019_015, w_015_089, w_017_004);
  and2 I019_016(w_019_016, w_013_158, w_004_138);
  nand2 I019_017(w_019_017, w_009_123, w_017_004);
  and2 I019_018(w_019_018, w_004_395, w_008_046);
  not1 I019_019(w_019_019, w_012_086);
  or2  I019_020(w_019_020, w_016_033, w_008_034);
  nand2 I019_021(w_019_021, w_008_020, w_017_025);
  or2  I019_022(w_019_022, w_015_129, w_013_123);
  nand2 I019_023(w_019_023, w_018_059, w_005_059);
  nand2 I019_024(w_019_024, w_003_053, w_007_055);
  and2 I019_025(w_019_025, w_012_358, w_011_077);
  and2 I019_026(w_019_026, w_017_179, w_014_034);
  or2  I019_027(w_019_027, w_017_071, w_011_213);
  or2  I019_028(w_019_028, w_013_194, w_017_188);
  nand2 I019_029(w_019_029, w_008_024, w_005_141);
  or2  I019_030(w_019_030, w_006_000, w_007_013);
  nand2 I019_031(w_019_031, w_003_088, w_013_017);
  nand2 I019_032(w_019_032, w_008_100, w_001_002);
  and2 I019_033(w_019_033, w_013_152, w_008_087);
  or2  I019_034(w_019_034, w_003_070, w_000_331);
  and2 I019_035(w_019_035, w_012_014, w_005_024);
  not1 I019_036(w_019_036, w_017_101);
  not1 I019_037(w_019_037, w_002_026);
  or2  I019_038(w_019_038, w_005_052, w_002_023);
  nand2 I019_039(w_019_039, w_007_180, w_011_020);
  and2 I019_040(w_019_040, w_006_000, w_009_010);
  not1 I019_041(w_019_041, w_009_034);
  not1 I019_042(w_019_042, w_011_246);
  or2  I019_043(w_019_043, w_017_099, w_002_005);
  or2  I019_044(w_019_044, w_016_303, w_006_000);
  and2 I019_045(w_019_045, w_009_148, w_010_219);
  not1 I019_046(w_019_046, w_017_059);
  nand2 I019_047(w_019_047, w_006_000, w_017_150);
  and2 I019_048(w_019_048, w_004_084, w_012_212);
  nand2 I019_049(w_019_049, w_004_459, w_001_006);
  not1 I019_050(w_019_050, w_000_346);
  and2 I019_051(w_019_051, w_017_001, w_007_083);
  not1 I019_052(w_019_052, w_016_374);
  or2  I019_053(w_019_053, w_002_004, w_011_096);
  nand2 I020_000(w_020_000, w_012_248, w_009_173);
  nand2 I020_001(w_020_001, w_005_055, w_011_304);
  nand2 I020_003(w_020_003, w_009_231, w_006_000);
  and2 I020_005(w_020_005, w_012_223, w_009_054);
  or2  I020_007(w_020_007, w_001_006, w_004_026);
  and2 I020_009(w_020_009, w_002_016, w_003_051);
  not1 I020_011(w_020_011, w_002_026);
  not1 I020_012(w_020_012, w_014_001);
  nand2 I020_013(w_020_013, w_007_194, w_005_050);
  not1 I020_014(w_020_014, w_007_128);
  nand2 I020_015(w_020_015, w_002_000, w_014_152);
  and2 I020_016(w_020_016, w_017_088, w_006_000);
  not1 I020_019(w_020_019, w_018_091);
  or2  I020_020(w_020_020, w_017_076, w_002_021);
  not1 I020_022(w_020_022, w_016_051);
  not1 I020_023(w_020_023, w_005_142);
  and2 I020_024(w_020_024, w_010_119, w_009_175);
  and2 I020_025(w_020_025, w_006_000, w_014_229);
  and2 I020_026(w_020_026, w_006_000, w_003_030);
  and2 I020_028(w_020_028, w_013_062, w_014_170);
  nand2 I020_030(w_020_030, w_015_115, w_018_016);
  not1 I020_031(w_020_031, w_002_010);
  not1 I020_032(w_020_032, w_016_079);
  nand2 I020_033(w_020_033, w_015_083, w_006_000);
  and2 I020_034(w_020_034, w_010_384, w_003_022);
  and2 I020_035(w_020_035, w_016_011, w_011_022);
  and2 I020_037(w_020_037, w_006_000, w_007_342);
  nand2 I020_038(w_020_038, w_009_096, w_006_000);
  nand2 I020_039(w_020_039, w_009_185, w_018_167);
  and2 I020_040(w_020_040, w_018_057, w_001_003);
  nand2 I020_042(w_020_042, w_012_166, w_016_023);
  or2  I020_043(w_020_043, w_017_157, w_010_336);
  nand2 I020_044(w_020_044, w_010_024, w_011_336);
  nand2 I020_045(w_020_045, w_003_081, w_012_221);
  and2 I020_046(w_020_046, w_001_000, w_001_005);
  and2 I020_048(w_020_048, w_019_012, w_016_324);
  not1 I020_049(w_020_049, w_012_347);
  nand2 I020_050(w_020_050, w_001_000, w_006_000);
  and2 I020_051(w_020_051, w_016_011, w_016_032);
  not1 I020_052(w_020_052, w_019_007);
  nand2 I020_053(w_020_053, w_012_090, w_008_184);
  not1 I020_054(w_020_054, w_002_010);
  or2  I020_055(w_020_055, w_013_122, w_005_244);
  nand2 I020_056(w_020_056, w_009_028, w_011_156);
  not1 I020_059(w_020_059, w_017_148);
  or2  I020_060(w_020_060, w_018_059, w_013_151);
  nand2 I020_062(w_020_062, w_002_011, w_016_152);
  not1 I020_063(w_020_063, w_005_180);
  nand2 I020_065(w_020_065, w_019_019, w_013_012);
  not1 I020_066(w_020_066, w_003_071);
  not1 I020_068(w_020_068, w_018_161);
  and2 I020_069(w_020_069, w_016_182, w_008_107);
  or2  I020_071(w_020_071, w_000_324, w_015_124);
  nand2 I020_072(w_020_072, w_007_305, w_013_268);
  nand2 I020_073(w_020_073, w_016_192, w_011_183);
  and2 I020_074(w_020_074, w_018_197, w_018_005);
  not1 I020_075(w_020_075, w_014_164);
  not1 I020_078(w_020_078, w_008_065);
  or2  I020_079(w_020_079, w_015_086, w_014_170);
  not1 I020_080(w_020_080, w_010_128);
  and2 I020_083(w_020_083, w_004_115, w_001_004);
  not1 I020_084(w_020_084, w_002_005);
  nand2 I020_085(w_020_085, w_015_067, w_004_421);
  and2 I020_086(w_020_086, w_011_143, w_007_007);
  and2 I020_088(w_020_088, w_010_309, w_015_042);
  not1 I020_089(w_020_089, w_004_021);
  nand2 I020_091(w_020_091, w_012_060, w_013_261);
  not1 I020_094(w_020_094, w_005_028);
  or2  I020_095(w_020_095, w_007_229, w_013_129);
  and2 I020_096(w_020_096, w_013_100, w_018_145);
  not1 I020_097(w_020_097, w_016_124);
  and2 I020_098(w_020_098, w_014_027, w_008_148);
  not1 I020_099(w_020_099, w_011_087);
  nand2 I020_100(w_020_100, w_002_024, w_016_228);
  not1 I020_101(w_020_101, w_017_042);
  or2  I020_103(w_020_103, w_005_047, w_002_001);
  or2  I020_104(w_020_104, w_002_020, w_013_046);
  and2 I020_105(w_020_105, w_007_192, w_008_133);
  not1 I020_106(w_020_106, w_012_221);
  or2  I020_107(w_020_107, w_014_195, w_017_030);
  and2 I020_108(w_020_108, w_006_000, w_000_263);
  and2 I020_112(w_020_112, w_002_024, w_018_074);
  or2  I020_113(w_020_113, w_000_260, w_018_257);
  not1 I020_114(w_020_114, w_002_016);
  nand2 I020_115(w_020_115, w_002_019, w_004_297);
  nand2 I020_117(w_020_117, w_004_436, w_012_215);
  not1 I020_119(w_020_119, w_016_026);
  nand2 I020_120(w_020_120, w_016_286, w_017_009);
  or2  I020_123(w_020_123, w_001_000, w_012_217);
  not1 I020_124(w_020_124, w_005_032);
  nand2 I020_125(w_020_125, w_015_031, w_004_195);
  or2  I020_126(w_020_126, w_000_221, w_012_328);
  nand2 I020_127(w_020_127, w_009_222, w_011_161);
  nand2 I020_128(w_020_128, w_003_004, w_004_280);
  not1 I020_131(w_020_131, w_009_208);
  and2 I020_135(w_020_135, w_012_373, w_009_046);
  or2  I020_136(w_020_136, w_000_095, w_015_052);
  nand2 I020_137(w_020_137, w_001_006, w_018_061);
  and2 I020_138(w_020_138, w_007_182, w_005_153);
  nand2 I020_139(w_020_139, w_008_086, w_013_174);
  nand2 I020_140(w_020_140, w_010_382, w_000_318);
  or2  I020_145(w_020_145, w_016_228, w_008_156);
  and2 I020_146(w_020_146, w_001_001, w_011_011);
  and2 I020_150(w_020_150, w_009_167, w_007_164);
  not1 I020_151(w_020_151, w_018_063);
  nand2 I020_152(w_020_152, w_006_000, w_011_215);
  not1 I020_153(w_020_153, w_004_398);
  or2  I020_154(w_020_154, w_007_058, w_004_408);
  or2  I020_155(w_020_155, w_016_264, w_000_365);
  nand2 I020_156(w_020_156, w_006_000, w_015_122);
  nand2 I020_157(w_020_157, w_016_061, w_014_206);
  nand2 I020_158(w_020_158, w_004_358, w_010_283);
  or2  I020_159(w_020_159, w_001_001, w_003_069);
  and2 I020_161(w_020_161, w_016_085, w_001_000);
  not1 I020_162(w_020_162, w_000_431);
  not1 I020_163(w_020_163, w_007_348);
  or2  I020_164(w_020_164, w_015_001, w_000_387);
  and2 I020_165(w_020_165, w_016_097, w_014_053);
  not1 I020_167(w_020_167, w_004_417);
  not1 I020_170(w_020_170, w_017_117);
  and2 I020_171(w_020_171, w_012_070, w_008_331);
  nand2 I020_172(w_020_172, w_004_428, w_001_000);
  nand2 I020_173(w_020_173, w_001_001, w_001_000);
  nand2 I020_175(w_020_175, w_017_018, w_005_003);
  nand2 I020_176(w_020_176, w_015_044, w_017_100);
  nand2 I020_180(w_020_180, w_003_092, w_018_108);
  not1 I020_182(w_020_182, w_012_068);
  or2  I020_183(w_020_183, w_007_119, w_015_051);
  and2 I020_184(w_020_184, w_000_139, w_016_254);
  not1 I020_186(w_020_186, w_014_144);
  nand2 I021_000(w_021_000, w_001_002, w_012_184);
  nand2 I021_001(w_021_001, w_018_282, w_020_127);
  not1 I021_002(w_021_002, w_016_106);
  not1 I021_003(w_021_003, w_005_014);
  or2  I021_005(w_021_005, w_009_203, w_002_000);
  not1 I021_007(w_021_007, w_012_322);
  and2 I021_008(w_021_008, w_013_245, w_006_000);
  or2  I021_009(w_021_009, w_003_039, w_006_000);
  nand2 I021_010(w_021_010, w_011_113, w_020_097);
  nand2 I021_011(w_021_011, w_004_432, w_003_075);
  or2  I021_012(w_021_012, w_003_069, w_020_094);
  or2  I021_014(w_021_014, w_002_002, w_014_066);
  or2  I021_015(w_021_015, w_004_059, w_000_002);
  nand2 I021_016(w_021_016, w_016_165, w_020_171);
  not1 I021_017(w_021_017, w_015_046);
  not1 I021_018(w_021_018, w_016_335);
  or2  I021_020(w_021_020, w_008_099, w_008_039);
  and2 I021_021(w_021_021, w_010_097, w_012_362);
  not1 I021_022(w_021_022, w_017_081);
  or2  I021_023(w_021_023, w_004_432, w_005_229);
  or2  I021_024(w_021_024, w_020_156, w_016_200);
  or2  I021_025(w_021_025, w_012_035, w_000_275);
  nand2 I021_026(w_021_026, w_019_047, w_005_191);
  not1 I021_027(w_021_027, w_013_231);
  not1 I021_028(w_021_028, w_001_006);
  and2 I021_029(w_021_029, w_016_247, w_012_171);
  and2 I021_030(w_021_030, w_017_072, w_011_276);
  or2  I021_031(w_021_031, w_008_120, w_015_013);
  or2  I021_032(w_021_032, w_006_000, w_008_130);
  nand2 I021_033(w_021_033, w_006_000, w_019_039);
  or2  I021_034(w_021_034, w_009_140, w_017_040);
  not1 I021_035(w_021_035, w_013_213);
  or2  I021_036(w_021_036, w_002_014, w_001_003);
  not1 I021_037(w_021_037, w_012_099);
  nand2 I021_038(w_021_038, w_020_080, w_016_034);
  nand2 I021_039(w_021_039, w_000_433, w_015_002);
  not1 I021_040(w_021_040, w_020_043);
  not1 I021_041(w_021_041, w_008_035);
  not1 I021_042(w_021_042, w_004_143);
  nand2 I021_043(w_021_043, w_005_171, w_007_386);
  or2  I021_044(w_021_044, w_007_023, w_012_070);
  and2 I021_045(w_021_045, w_006_000, w_012_088);
  and2 I021_047(w_021_047, w_013_211, w_005_222);
  not1 I021_048(w_021_048, w_013_094);
  or2  I021_049(w_021_049, w_017_006, w_003_051);
  or2  I021_050(w_021_050, w_008_345, w_001_004);
  or2  I021_051(w_021_051, w_013_110, w_014_262);
  nand2 I021_052(w_021_052, w_003_029, w_005_189);
  and2 I021_053(w_021_053, w_005_065, w_020_040);
  and2 I021_056(w_021_056, w_019_036, w_005_075);
  nand2 I021_057(w_021_057, w_006_000, w_002_008);
  and2 I021_058(w_021_058, w_007_074, w_010_153);
  or2  I021_059(w_021_059, w_001_006, w_011_151);
  and2 I021_060(w_021_060, w_007_058, w_013_227);
  or2  I021_061(w_021_061, w_010_096, w_020_062);
  nand2 I021_063(w_021_063, w_005_130, w_010_433);
  nand2 I021_064(w_021_064, w_017_058, w_010_067);
  nand2 I021_066(w_021_066, w_004_316, w_001_006);
  and2 I021_067(w_021_067, w_014_156, w_013_148);
  and2 I021_069(w_021_069, w_001_001, w_019_019);
  nand2 I021_070(w_021_070, w_009_096, w_003_013);
  and2 I021_071(w_021_071, w_001_001, w_011_092);
  or2  I021_072(w_021_072, w_013_071, w_016_107);
  or2  I021_073(w_021_073, w_019_015, w_019_044);
  not1 I021_075(w_021_075, w_018_150);
  and2 I021_076(w_021_076, w_016_101, w_000_032);
  not1 I021_077(w_021_077, w_001_005);
  not1 I021_078(w_021_078, w_002_026);
  nand2 I021_079(w_021_079, w_018_200, w_010_270);
  and2 I021_081(w_021_081, w_008_138, w_014_207);
  not1 I021_082(w_021_082, w_008_196);
  not1 I021_083(w_021_083, w_006_000);
  or2  I021_084(w_021_084, w_013_049, w_017_044);
  not1 I021_085(w_021_085, w_014_227);
  and2 I021_086(w_021_086, w_000_330, w_018_047);
  not1 I021_088(w_021_088, w_009_145);
  or2  I021_089(w_021_089, w_013_083, w_015_077);
  not1 I021_090(w_021_090, w_010_034);
  and2 I021_091(w_021_091, w_002_016, w_013_060);
  nand2 I021_092(w_021_092, w_006_000, w_001_001);
  nand2 I021_093(w_021_093, w_000_069, w_019_038);
  not1 I021_094(w_021_094, w_003_006);
  not1 I021_096(w_021_096, w_006_000);
  nand2 I021_097(w_021_097, w_004_097, w_017_003);
  or2  I021_098(w_021_098, w_017_187, w_003_006);
  not1 I021_099(w_021_099, w_007_325);
  not1 I021_100(w_021_100, w_005_096);
  and2 I021_101(w_021_101, w_017_018, w_013_007);
  nand2 I021_102(w_021_102, w_011_220, w_015_059);
  nand2 I021_103(w_021_103, w_003_002, w_019_046);
  or2  I021_104(w_021_104, w_002_019, w_007_344);
  and2 I021_105(w_021_105, w_003_076, w_017_087);
  not1 I021_106(w_021_106, w_003_048);
  and2 I021_107(w_021_107, w_007_404, w_000_040);
  not1 I021_108(w_021_108, w_011_047);
  or2  I021_109(w_021_109, w_000_119, w_002_022);
  not1 I022_000(w_022_000, w_014_216);
  or2  I022_002(w_022_002, w_019_033, w_009_026);
  nand2 I022_003(w_022_003, w_000_066, w_021_102);
  or2  I022_004(w_022_004, w_004_018, w_016_048);
  and2 I022_005(w_022_005, w_002_006, w_000_315);
  nand2 I022_006(w_022_006, w_008_241, w_021_090);
  nand2 I022_007(w_022_007, w_011_031, w_006_000);
  not1 I022_009(w_022_009, w_000_196);
  or2  I022_010(w_022_010, w_000_114, w_021_097);
  nand2 I022_011(w_022_011, w_003_064, w_011_035);
  not1 I022_012(w_022_012, w_013_135);
  nand2 I022_013(w_022_013, w_010_063, w_019_053);
  not1 I022_014(w_022_014, w_016_133);
  or2  I022_016(w_022_016, w_001_003, w_021_015);
  or2  I022_018(w_022_018, w_009_030, w_012_180);
  and2 I022_020(w_022_020, w_020_138, w_015_091);
  nand2 I022_021(w_022_021, w_004_458, w_005_191);
  and2 I022_023(w_022_023, w_016_191, w_015_063);
  and2 I022_024(w_022_024, w_014_164, w_006_000);
  and2 I022_025(w_022_025, w_000_122, w_019_035);
  or2  I022_027(w_022_027, w_005_246, w_013_165);
  not1 I022_028(w_022_028, w_005_105);
  or2  I022_032(w_022_032, w_000_085, w_012_110);
  not1 I022_033(w_022_033, w_004_286);
  nand2 I022_034(w_022_034, w_007_285, w_018_012);
  nand2 I022_035(w_022_035, w_001_005, w_008_013);
  or2  I022_036(w_022_036, w_018_133, w_000_342);
  and2 I022_037(w_022_037, w_021_099, w_011_140);
  or2  I022_038(w_022_038, w_014_222, w_000_434);
  and2 I022_040(w_022_040, w_013_088, w_019_033);
  nand2 I022_041(w_022_041, w_010_315, w_004_217);
  and2 I022_042(w_022_042, w_017_171, w_014_235);
  or2  I022_043(w_022_043, w_002_010, w_004_406);
  nand2 I022_044(w_022_044, w_014_106, w_019_028);
  and2 I022_046(w_022_046, w_017_018, w_012_000);
  or2  I022_049(w_022_049, w_000_096, w_009_088);
  not1 I022_050(w_022_050, w_002_012);
  not1 I022_051(w_022_051, w_021_109);
  nand2 I022_052(w_022_052, w_017_150, w_006_000);
  nand2 I022_053(w_022_053, w_021_103, w_011_017);
  nand2 I022_055(w_022_055, w_004_473, w_016_291);
  not1 I022_056(w_022_056, w_016_239);
  or2  I022_057(w_022_057, w_016_093, w_006_000);
  and2 I022_058(w_022_058, w_003_054, w_017_047);
  and2 I022_059(w_022_059, w_002_004, w_015_043);
  nand2 I022_062(w_022_062, w_020_071, w_011_228);
  and2 I022_064(w_022_064, w_018_106, w_008_152);
  and2 I022_065(w_022_065, w_003_083, w_018_237);
  not1 I022_067(w_022_067, w_005_245);
  not1 I022_069(w_022_069, w_014_129);
  nand2 I022_070(w_022_070, w_004_292, w_002_011);
  and2 I022_071(w_022_071, w_020_042, w_020_034);
  or2  I022_072(w_022_072, w_021_007, w_018_010);
  or2  I022_074(w_022_074, w_019_038, w_020_091);
  or2  I022_075(w_022_075, w_019_002, w_000_420);
  and2 I022_076(w_022_076, w_014_049, w_020_162);
  not1 I022_078(w_022_078, w_003_027);
  nand2 I022_079(w_022_079, w_003_074, w_001_006);
  and2 I022_081(w_022_081, w_018_291, w_009_080);
  or2  I022_082(w_022_082, w_007_090, w_003_056);
  nand2 I022_083(w_022_083, w_001_004, w_013_046);
  or2  I022_084(w_022_084, w_020_007, w_005_059);
  or2  I022_085(w_022_085, w_009_089, w_005_044);
  or2  I022_088(w_022_088, w_010_004, w_001_000);
  nand2 I022_090(w_022_090, w_000_422, w_011_016);
  not1 I022_091(w_022_091, w_004_402);
  nand2 I022_092(w_022_092, w_009_209, w_018_142);
  nand2 I022_093(w_022_093, w_011_336, w_003_058);
  or2  I022_095(w_022_095, w_017_101, w_007_066);
  or2  I022_096(w_022_096, w_007_005, w_004_117);
  nand2 I022_098(w_022_098, w_004_448, w_000_266);
  not1 I022_099(w_022_099, w_013_267);
  nand2 I022_101(w_022_101, w_015_111, w_017_182);
  or2  I022_102(w_022_102, w_002_024, w_014_087);
  not1 I022_103(w_022_103, w_016_067);
  nand2 I022_105(w_022_105, w_007_045, w_004_058);
  or2  I022_106(w_022_106, w_015_053, w_018_072);
  or2  I022_107(w_022_107, w_016_068, w_000_105);
  and2 I022_109(w_022_109, w_017_167, w_002_001);
  not1 I022_110(w_022_110, w_012_312);
  or2  I022_112(w_022_112, w_002_012, w_021_052);
  or2  I022_113(w_022_113, w_015_046, w_013_046);
  nand2 I022_114(w_022_114, w_008_288, w_019_009);
  and2 I022_115(w_022_115, w_013_096, w_009_080);
  not1 I022_116(w_022_116, w_004_010);
  and2 I022_117(w_022_117, w_013_123, w_000_289);
  or2  I022_118(w_022_118, w_015_047, w_015_002);
  and2 I022_120(w_022_120, w_008_121, w_017_030);
  or2  I022_121(w_022_121, w_015_120, w_015_072);
  or2  I022_122(w_022_122, w_002_026, w_005_177);
  and2 I022_123(w_022_123, w_014_141, w_019_024);
  and2 I022_124(w_022_124, w_013_012, w_001_000);
  and2 I022_126(w_022_126, w_013_099, w_021_102);
  or2  I022_127(w_022_127, w_014_096, w_018_168);
  or2  I022_131(w_022_131, w_020_020, w_000_406);
  or2  I022_132(w_022_132, w_004_396, w_021_101);
  and2 I022_133(w_022_133, w_013_164, w_021_041);
  not1 I022_134(w_022_134, w_014_085);
  or2  I022_137(w_022_137, w_013_177, w_002_017);
  nand2 I022_138(w_022_138, w_001_006, w_014_043);
  nand2 I022_139(w_022_139, w_011_108, w_015_078);
  or2  I022_140(w_022_140, w_013_055, w_007_315);
  or2  I022_141(w_022_141, w_007_324, w_007_021);
  or2  I022_142(w_022_142, w_015_046, w_002_004);
  or2  I022_143(w_022_143, w_015_047, w_006_000);
  and2 I022_144(w_022_144, w_017_041, w_011_078);
  and2 I022_145(w_022_145, w_002_025, w_001_005);
  nand2 I022_146(w_022_146, w_002_019, w_005_193);
  not1 I022_147(w_022_147, w_014_137);
  not1 I022_148(w_022_148, w_019_010);
  and2 I022_149(w_022_149, w_012_234, w_008_098);
  not1 I022_152(w_022_152, w_003_059);
  nand2 I022_154(w_022_154, w_007_008, w_017_091);
  not1 I022_156(w_022_156, w_020_161);
  not1 I022_157(w_022_157, w_006_000);
  and2 I022_158(w_022_158, w_004_311, w_002_013);
  nand2 I022_159(w_022_159, w_011_112, w_007_261);
  nand2 I022_160(w_022_160, w_005_156, w_014_049);
  and2 I022_161(w_022_161, w_019_044, w_005_047);
  nand2 I022_162(w_022_162, w_014_109, w_009_112);
  or2  I022_163(w_022_165, w_002_020, w_022_164);
  and2 I022_164(w_022_166, w_022_165, w_010_284);
  and2 I022_165(w_022_167, w_022_166, w_018_060);
  or2  I022_166(w_022_168, w_022_167, w_018_295);
  nand2 I022_167(w_022_169, w_011_219, w_022_168);
  nand2 I022_168(w_022_170, w_004_034, w_022_169);
  nand2 I022_169(w_022_171, w_022_170, w_004_360);
  or2  I022_170(w_022_172, w_021_107, w_022_171);
  and2 I022_171(w_022_173, w_014_264, w_022_172);
  or2  I022_172(w_022_164, w_012_197, w_022_173);
  or2  I023_000(w_023_000, w_002_025, w_006_000);
  and2 I023_002(w_023_002, w_004_455, w_021_020);
  not1 I023_006(w_023_006, w_009_075);
  nand2 I023_009(w_023_009, w_017_012, w_009_132);
  not1 I023_010(w_023_010, w_020_035);
  not1 I023_013(w_023_013, w_002_001);
  not1 I023_014(w_023_014, w_004_430);
  or2  I023_016(w_023_016, w_004_350, w_010_042);
  and2 I023_018(w_023_018, w_010_069, w_007_078);
  nand2 I023_020(w_023_020, w_001_003, w_020_013);
  not1 I023_024(w_023_024, w_003_039);
  not1 I023_028(w_023_028, w_015_012);
  nand2 I023_030(w_023_030, w_012_094, w_016_124);
  or2  I023_031(w_023_031, w_003_085, w_010_127);
  and2 I023_034(w_023_034, w_012_046, w_022_088);
  not1 I023_038(w_023_038, w_020_120);
  nand2 I023_039(w_023_039, w_009_009, w_019_025);
  not1 I023_041(w_023_041, w_015_021);
  and2 I023_042(w_023_042, w_016_194, w_022_156);
  or2  I023_043(w_023_043, w_011_022, w_009_132);
  and2 I023_046(w_023_046, w_004_168, w_020_135);
  or2  I023_047(w_023_047, w_000_258, w_013_225);
  and2 I023_049(w_023_049, w_016_176, w_004_011);
  and2 I023_050(w_023_050, w_010_152, w_005_074);
  not1 I023_051(w_023_051, w_017_108);
  nand2 I023_052(w_023_052, w_002_026, w_014_220);
  not1 I023_053(w_023_053, w_006_000);
  or2  I023_058(w_023_058, w_018_155, w_022_093);
  not1 I023_059(w_023_059, w_008_130);
  or2  I023_061(w_023_061, w_002_024, w_003_035);
  nand2 I023_063(w_023_063, w_021_022, w_018_213);
  not1 I023_064(w_023_064, w_002_000);
  not1 I023_067(w_023_067, w_020_158);
  nand2 I023_068(w_023_068, w_022_160, w_009_217);
  not1 I023_071(w_023_071, w_002_007);
  nand2 I023_072(w_023_072, w_009_117, w_000_437);
  or2  I023_074(w_023_074, w_022_105, w_022_156);
  nand2 I023_075(w_023_075, w_021_031, w_000_155);
  not1 I023_081(w_023_081, w_000_431);
  or2  I023_082(w_023_082, w_015_126, w_022_078);
  and2 I023_083(w_023_083, w_001_005, w_018_302);
  nand2 I023_100(w_023_100, w_020_030, w_004_167);
  not1 I023_104(w_023_104, w_005_058);
  not1 I023_110(w_023_110, w_007_270);
  not1 I023_120(w_023_120, w_022_056);
  not1 I023_121(w_023_121, w_008_082);
  nand2 I023_122(w_023_122, w_004_023, w_003_022);
  or2  I023_126(w_023_126, w_009_064, w_019_032);
  nand2 I023_137(w_023_137, w_003_071, w_018_314);
  nand2 I023_138(w_023_138, w_005_021, w_020_050);
  and2 I023_140(w_023_140, w_007_039, w_013_027);
  nand2 I023_144(w_023_144, w_001_006, w_018_215);
  and2 I023_145(w_023_145, w_020_107, w_002_004);
  nand2 I023_150(w_023_150, w_002_026, w_001_000);
  or2  I023_156(w_023_156, w_009_007, w_008_187);
  and2 I023_159(w_023_159, w_019_022, w_018_162);
  nand2 I023_161(w_023_161, w_014_001, w_018_026);
  or2  I023_163(w_023_163, w_011_028, w_007_231);
  not1 I023_165(w_023_165, w_008_092);
  or2  I023_172(w_023_172, w_018_302, w_005_237);
  not1 I023_176(w_023_176, w_017_114);
  or2  I023_177(w_023_177, w_000_004, w_003_092);
  nand2 I023_179(w_023_179, w_003_061, w_007_288);
  nand2 I023_180(w_023_180, w_021_010, w_019_003);
  or2  I023_182(w_023_182, w_016_058, w_021_108);
  and2 I023_183(w_023_183, w_016_058, w_017_088);
  and2 I023_185(w_023_185, w_022_065, w_015_075);
  and2 I023_189(w_023_189, w_014_088, w_016_080);
  and2 I023_190(w_023_190, w_011_116, w_001_004);
  not1 I023_191(w_023_191, w_014_040);
  not1 I023_192(w_023_192, w_007_063);
  or2  I023_196(w_023_196, w_018_032, w_006_000);
  or2  I023_197(w_023_197, w_017_081, w_010_315);
  and2 I023_201(w_023_201, w_004_316, w_014_198);
  nand2 I023_209(w_023_209, w_011_268, w_002_019);
  and2 I023_210(w_023_210, w_011_057, w_011_043);
  and2 I023_215(w_023_215, w_001_002, w_000_257);
  or2  I023_218(w_023_218, w_007_117, w_021_093);
  and2 I023_220(w_023_220, w_000_413, w_004_135);
  and2 I023_228(w_023_228, w_015_122, w_014_110);
  not1 I023_231(w_023_231, w_012_169);
  or2  I023_232(w_023_232, w_001_003, w_006_000);
  and2 I023_233(w_023_233, w_021_049, w_019_037);
  and2 I023_235(w_023_235, w_005_217, w_013_059);
  nand2 I023_238(w_023_238, w_007_082, w_017_034);
  or2  I023_239(w_023_239, w_016_058, w_016_091);
  or2  I023_244(w_023_244, w_003_008, w_019_022);
  nand2 I023_251(w_023_251, w_006_000, w_010_181);
  nand2 I023_256(w_023_256, w_015_096, w_014_118);
  nand2 I023_259(w_023_259, w_005_137, w_005_059);
  not1 I023_264(w_023_264, w_009_007);
  or2  I023_267(w_023_267, w_002_016, w_001_001);
  or2  I023_269(w_023_269, w_008_270, w_005_032);
  not1 I023_270(w_023_270, w_000_368);
  and2 I023_271(w_023_271, w_009_204, w_001_002);
  and2 I023_272(w_023_272, w_002_007, w_020_095);
  nand2 I023_275(w_023_275, w_019_004, w_021_089);
  not1 I023_277(w_023_277, w_013_171);
  and2 I023_284(w_023_284, w_018_089, w_014_008);
  not1 I023_285(w_023_285, w_016_101);
  nand2 I023_290(w_023_290, w_011_076, w_010_185);
  and2 I023_295(w_023_295, w_006_000, w_010_142);
  nand2 I023_301(w_023_301, w_004_341, w_012_182);
  not1 I023_306(w_023_306, w_004_421);
  not1 I023_307(w_023_307, w_009_193);
  nand2 I023_309(w_023_309, w_018_008, w_018_060);
  and2 I023_311(w_023_311, w_016_031, w_009_086);
  or2  I023_312(w_023_312, w_010_278, w_004_143);
  not1 I023_314(w_023_314, w_017_040);
  and2 I023_318(w_023_318, w_016_026, w_022_023);
  nand2 I023_319(w_023_319, w_010_026, w_001_005);
  nand2 I023_323(w_023_323, w_007_307, w_010_303);
  nand2 I023_324(w_023_324, w_001_006, w_006_000);
  or2  I023_325(w_023_325, w_009_171, w_011_156);
  nand2 I023_327(w_023_327, w_016_007, w_013_059);
  nand2 I023_330(w_023_330, w_020_117, w_022_157);
  or2  I023_334(w_023_334, w_002_015, w_000_312);
  and2 I023_335(w_023_335, w_005_053, w_014_076);
  and2 I023_340(w_023_340, w_020_033, w_005_087);
  or2  I023_348(w_023_348, w_003_088, w_017_014);
  nand2 I023_350(w_023_350, w_006_000, w_015_117);
  not1 I023_351(w_023_351, w_003_046);
  nand2 I023_353(w_023_353, w_001_000, w_018_133);
  nand2 I023_354(w_023_354, w_007_241, w_000_061);
  nand2 I023_359(w_023_359, w_011_233, w_002_020);
  nand2 I023_367(w_023_367, w_015_077, w_001_002);
  and2 I023_369(w_023_369, w_003_044, w_001_002);
  and2 I023_373(w_023_373, w_014_027, w_008_070);
  nand2 I023_374(w_023_374, w_020_011, w_022_140);
  or2  I023_376(w_023_376, w_006_000, w_001_005);
  or2  I023_379(w_023_379, w_014_207, w_021_083);
  not1 I023_386(w_023_386, w_019_033);
  nand2 I023_388(w_023_388, w_009_014, w_006_000);
  not1 I023_393(w_023_393, w_012_149);
  and2 I023_395(w_023_395, w_017_053, w_000_440);
  and2 I023_400(w_023_400, w_009_226, w_015_045);
  or2  I023_401(w_023_401, w_018_114, w_001_001);
  nand2 I023_402(w_023_402, w_018_313, w_002_027);
  nand2 I023_404(w_023_404, w_008_105, w_022_055);
  nand2 I023_413(w_023_413, w_013_024, w_003_001);
  or2  I024_000(w_024_000, w_014_074, w_010_120);
  nand2 I024_002(w_024_002, w_004_441, w_005_100);
  and2 I024_003(w_024_003, w_005_014, w_019_047);
  not1 I024_004(w_024_004, w_011_120);
  nand2 I024_007(w_024_007, w_015_007, w_011_077);
  or2  I024_008(w_024_008, w_009_206, w_005_032);
  and2 I024_009(w_024_009, w_010_385, w_012_043);
  or2  I024_016(w_024_016, w_017_178, w_013_011);
  or2  I024_018(w_024_018, w_003_010, w_022_113);
  nand2 I024_019(w_024_019, w_009_154, w_002_012);
  or2  I024_021(w_024_021, w_018_134, w_005_113);
  and2 I024_023(w_024_023, w_011_000, w_011_166);
  not1 I024_025(w_024_025, w_010_380);
  nand2 I024_027(w_024_027, w_017_091, w_021_067);
  nand2 I024_031(w_024_031, w_017_117, w_019_020);
  nand2 I024_032(w_024_032, w_005_000, w_019_000);
  not1 I024_033(w_024_033, w_014_070);
  or2  I024_036(w_024_036, w_016_232, w_006_000);
  not1 I024_037(w_024_037, w_018_211);
  not1 I024_040(w_024_040, w_005_170);
  nand2 I024_042(w_024_042, w_015_017, w_004_187);
  not1 I024_044(w_024_044, w_000_254);
  and2 I024_045(w_024_045, w_004_136, w_012_320);
  or2  I024_046(w_024_046, w_021_072, w_015_054);
  nand2 I024_048(w_024_048, w_014_053, w_016_279);
  not1 I024_049(w_024_049, w_007_148);
  and2 I024_051(w_024_051, w_009_134, w_021_027);
  and2 I024_052(w_024_052, w_001_001, w_013_061);
  and2 I024_053(w_024_053, w_010_321, w_020_005);
  and2 I024_054(w_024_054, w_008_294, w_007_226);
  or2  I024_055(w_024_055, w_015_085, w_004_418);
  not1 I024_057(w_024_057, w_005_198);
  nand2 I024_058(w_024_058, w_014_156, w_012_318);
  nand2 I024_059(w_024_059, w_005_169, w_016_322);
  not1 I024_060(w_024_060, w_018_173);
  not1 I024_061(w_024_061, w_010_368);
  or2  I024_064(w_024_064, w_012_373, w_002_011);
  not1 I024_065(w_024_065, w_012_003);
  or2  I024_066(w_024_066, w_007_001, w_003_030);
  nand2 I024_067(w_024_067, w_000_222, w_017_042);
  and2 I024_068(w_024_068, w_017_028, w_014_205);
  nand2 I024_069(w_024_069, w_015_073, w_012_270);
  and2 I024_070(w_024_070, w_022_162, w_021_007);
  not1 I024_071(w_024_071, w_015_050);
  and2 I024_072(w_024_072, w_020_157, w_013_267);
  not1 I024_073(w_024_073, w_008_205);
  or2  I024_074(w_024_074, w_001_006, w_018_156);
  nand2 I024_075(w_024_075, w_012_052, w_001_006);
  nand2 I024_076(w_024_076, w_009_134, w_015_063);
  and2 I024_078(w_024_078, w_016_265, w_003_004);
  or2  I024_081(w_024_081, w_005_070, w_008_228);
  not1 I024_084(w_024_084, w_020_123);
  not1 I024_085(w_024_085, w_004_428);
  not1 I024_086(w_024_086, w_023_126);
  or2  I024_087(w_024_087, w_017_077, w_016_078);
  or2  I024_088(w_024_088, w_015_047, w_002_002);
  nand2 I024_089(w_024_089, w_019_003, w_023_179);
  not1 I024_090(w_024_090, w_021_027);
  not1 I024_093(w_024_093, w_000_068);
  nand2 I024_096(w_024_096, w_023_163, w_018_094);
  not1 I024_100(w_024_100, w_003_075);
  or2  I024_103(w_024_103, w_017_076, w_020_025);
  nand2 I024_105(w_024_105, w_001_004, w_003_038);
  and2 I024_106(w_024_106, w_017_059, w_003_066);
  or2  I024_109(w_024_109, w_007_296, w_019_005);
  and2 I024_110(w_024_110, w_007_364, w_001_003);
  or2  I024_111(w_024_111, w_006_000, w_004_295);
  nand2 I024_112(w_024_112, w_007_038, w_000_288);
  or2  I024_114(w_024_114, w_009_018, w_005_049);
  or2  I024_115(w_024_115, w_014_145, w_010_265);
  not1 I024_116(w_024_116, w_014_209);
  not1 I024_117(w_024_117, w_016_345);
  or2  I024_121(w_024_121, w_022_037, w_007_276);
  not1 I024_122(w_024_122, w_013_153);
  nand2 I024_123(w_024_123, w_007_007, w_016_249);
  or2  I024_124(w_024_124, w_010_283, w_006_000);
  or2  I024_127(w_024_127, w_009_179, w_014_193);
  and2 I024_128(w_024_128, w_013_235, w_006_000);
  nand2 I024_130(w_024_130, w_005_052, w_018_032);
  not1 I024_131(w_024_131, w_002_006);
  not1 I024_132(w_024_132, w_023_351);
  not1 I024_133(w_024_133, w_010_379);
  nand2 I024_135(w_024_135, w_021_105, w_008_329);
  nand2 I024_136(w_024_136, w_003_069, w_009_233);
  or2  I024_139(w_024_139, w_012_048, w_012_367);
  not1 I024_140(w_024_140, w_001_000);
  or2  I024_143(w_024_143, w_017_187, w_022_152);
  and2 I024_144(w_024_144, w_014_221, w_003_015);
  nand2 I024_148(w_024_148, w_020_119, w_021_084);
  or2  I024_150(w_024_150, w_020_108, w_001_006);
  nand2 I024_151(w_024_151, w_020_020, w_005_036);
  or2  I024_152(w_024_152, w_013_180, w_005_008);
  and2 I024_153(w_024_153, w_009_020, w_009_004);
  not1 I024_163(w_024_163, w_003_035);
  not1 I024_164(w_024_164, w_014_040);
  not1 I024_165(w_024_165, w_021_088);
  nand2 I024_166(w_024_166, w_014_184, w_009_125);
  not1 I024_169(w_024_169, w_023_393);
  nand2 I024_170(w_024_170, w_004_233, w_012_023);
  or2  I024_173(w_024_173, w_010_047, w_022_055);
  or2  I024_174(w_024_174, w_014_037, w_018_197);
  or2  I024_176(w_024_176, w_014_260, w_008_251);
  or2  I024_177(w_024_177, w_020_009, w_012_110);
  not1 I024_178(w_024_178, w_015_014);
  or2  I024_179(w_024_179, w_022_159, w_021_025);
  not1 I024_180(w_024_180, w_008_260);
  or2  I024_181(w_024_181, w_006_000, w_011_114);
  and2 I024_182(w_024_182, w_021_063, w_019_009);
  and2 I024_183(w_024_183, w_009_147, w_016_152);
  nand2 I024_185(w_024_185, w_012_133, w_016_110);
  not1 I024_186(w_024_186, w_014_057);
  and2 I024_187(w_024_187, w_014_084, w_005_152);
  not1 I024_188(w_024_188, w_017_077);
  not1 I024_189(w_024_189, w_014_024);
  or2  I024_190(w_024_190, w_017_065, w_010_009);
  or2  I024_191(w_024_191, w_007_354, w_022_137);
  and2 I024_194(w_024_194, w_000_226, w_017_064);
  not1 I024_196(w_024_196, w_011_126);
  nand2 I024_197(w_024_197, w_021_039, w_004_112);
  nand2 I024_205(w_024_205, w_023_197, w_004_095);
  not1 I024_206(w_024_206, w_013_150);
  nand2 I024_209(w_024_209, w_015_041, w_015_093);
  not1 I024_210(w_024_210, w_000_118);
  not1 I024_211(w_024_211, w_002_021);
  or2  I024_214(w_024_214, w_007_025, w_007_309);
  nand2 I024_216(w_024_216, w_005_134, w_022_083);
  or2  I024_217(w_024_217, w_014_216, w_012_021);
  not1 I024_222(w_024_222, w_020_051);
  not1 I024_226(w_024_226, w_023_386);
  not1 I024_228(w_024_228, w_015_066);
  nand2 I024_229(w_024_229, w_014_067, w_001_005);
  and2 I024_230(w_024_230, w_002_009, w_006_000);
  not1 I024_235(w_024_235, w_000_023);
  or2  I024_239(w_024_239, w_020_037, w_007_082);
  and2 I024_240(w_024_240, w_014_157, w_004_076);
  nand2 I024_241(w_024_241, w_011_342, w_018_070);
  not1 I024_244(w_024_244, w_011_205);
  nand2 I024_245(w_024_245, w_013_019, w_004_313);
  not1 I024_249(w_024_249, w_001_001);
  or2  I024_250(w_024_250, w_000_381, w_015_074);
  and2 I024_251(w_024_251, w_002_023, w_015_048);
  and2 I024_258(w_024_258, w_002_016, w_003_074);
  not1 I024_259(w_024_259, w_014_115);
  and2 I024_261(w_024_261, w_015_077, w_021_056);
  nand2 I024_266(w_024_266, w_009_084, w_008_032);
  not1 I024_270(w_024_270, w_003_087);
  nand2 I024_275(w_024_275, w_020_158, w_021_082);
  and2 I024_276(w_024_276, w_005_188, w_004_102);
  not1 I024_277(w_024_277, w_023_144);
  and2 I024_280(w_024_280, w_021_049, w_019_027);
  not1 I024_284(w_024_284, w_019_013);
  and2 I024_285(w_024_285, w_013_221, w_007_246);
  not1 I024_287(w_024_287, w_012_023);
  nand2 I024_294(w_024_294, w_011_085, w_008_015);
  nand2 I024_295(w_024_295, w_004_444, w_018_027);
  not1 I024_296(w_024_296, w_019_047);
  or2  I024_297(w_024_297, w_002_010, w_014_133);
  nand2 I025_007(w_025_007, w_021_044, w_008_089);
  nand2 I025_009(w_025_009, w_010_413, w_008_096);
  not1 I025_010(w_025_010, w_005_199);
  nand2 I025_012(w_025_012, w_023_042, w_016_062);
  nand2 I025_013(w_025_013, w_001_004, w_008_299);
  not1 I025_014(w_025_014, w_017_004);
  or2  I025_015(w_025_015, w_012_283, w_019_048);
  not1 I025_016(w_025_016, w_005_069);
  nand2 I025_017(w_025_017, w_001_001, w_000_354);
  and2 I025_019(w_025_019, w_016_094, w_010_234);
  or2  I025_020(w_025_020, w_013_159, w_002_005);
  nand2 I025_023(w_025_023, w_011_312, w_018_040);
  not1 I025_026(w_025_026, w_001_001);
  or2  I025_029(w_025_029, w_012_171, w_018_279);
  not1 I025_030(w_025_030, w_007_038);
  not1 I025_045(w_025_045, w_009_159);
  not1 I025_056(w_025_056, w_012_175);
  and2 I025_060(w_025_060, w_000_151, w_021_039);
  not1 I025_063(w_025_063, w_023_067);
  not1 I025_066(w_025_066, w_020_097);
  or2  I025_069(w_025_069, w_020_044, w_010_132);
  nand2 I025_070(w_025_070, w_000_118, w_000_278);
  not1 I025_071(w_025_071, w_017_187);
  not1 I025_073(w_025_073, w_019_033);
  and2 I025_074(w_025_074, w_016_086, w_009_111);
  not1 I025_079(w_025_079, w_017_063);
  not1 I025_082(w_025_082, w_024_217);
  and2 I025_085(w_025_085, w_012_092, w_020_151);
  nand2 I025_089(w_025_089, w_010_059, w_001_004);
  not1 I025_091(w_025_091, w_001_001);
  nand2 I025_092(w_025_092, w_013_081, w_003_061);
  nand2 I025_093(w_025_093, w_021_003, w_015_089);
  not1 I025_094(w_025_094, w_008_123);
  not1 I025_095(w_025_095, w_006_000);
  and2 I025_097(w_025_097, w_017_012, w_019_014);
  not1 I025_101(w_025_101, w_015_000);
  nand2 I025_104(w_025_104, w_005_026, w_023_064);
  not1 I025_105(w_025_105, w_004_460);
  not1 I025_106(w_025_106, w_018_063);
  and2 I025_113(w_025_113, w_004_440, w_015_005);
  or2  I025_115(w_025_115, w_001_000, w_015_069);
  and2 I025_127(w_025_127, w_024_297, w_006_000);
  not1 I025_130(w_025_130, w_007_321);
  nand2 I025_137(w_025_137, w_002_024, w_001_006);
  or2  I025_143(w_025_143, w_024_239, w_020_125);
  and2 I025_146(w_025_146, w_018_104, w_023_259);
  or2  I025_149(w_025_149, w_013_039, w_012_362);
  not1 I025_150(w_025_150, w_007_174);
  and2 I025_155(w_025_155, w_011_093, w_008_246);
  not1 I025_156(w_025_156, w_023_137);
  nand2 I025_159(w_025_159, w_020_128, w_005_151);
  not1 I025_160(w_025_160, w_006_000);
  not1 I025_165(w_025_165, w_015_026);
  or2  I025_172(w_025_172, w_008_277, w_007_122);
  or2  I025_174(w_025_174, w_008_186, w_014_059);
  and2 I025_180(w_025_180, w_022_147, w_002_017);
  nand2 I025_190(w_025_190, w_007_225, w_013_024);
  nand2 I025_194(w_025_194, w_013_104, w_010_008);
  nand2 I025_195(w_025_195, w_004_285, w_008_302);
  and2 I025_197(w_025_197, w_011_315, w_006_000);
  or2  I025_200(w_025_200, w_002_023, w_017_080);
  not1 I025_212(w_025_212, w_010_023);
  and2 I025_214(w_025_214, w_009_042, w_000_378);
  or2  I025_220(w_025_220, w_006_000, w_003_004);
  and2 I025_226(w_025_226, w_002_023, w_006_000);
  not1 I025_233(w_025_233, w_007_374);
  nand2 I025_234(w_025_234, w_014_035, w_013_030);
  nand2 I025_237(w_025_237, w_017_010, w_004_314);
  nand2 I025_240(w_025_240, w_017_064, w_018_182);
  or2  I025_244(w_025_244, w_003_044, w_009_098);
  and2 I025_245(w_025_245, w_016_250, w_021_069);
  or2  I025_248(w_025_248, w_006_000, w_010_123);
  nand2 I025_249(w_025_249, w_013_207, w_006_000);
  not1 I025_258(w_025_258, w_017_146);
  nand2 I025_260(w_025_260, w_015_004, w_017_066);
  or2  I025_261(w_025_261, w_013_152, w_019_025);
  not1 I025_262(w_025_262, w_003_081);
  not1 I025_264(w_025_264, w_011_323);
  or2  I025_265(w_025_265, w_019_041, w_007_341);
  nand2 I025_275(w_025_275, w_021_034, w_015_071);
  not1 I025_276(w_025_276, w_023_201);
  not1 I025_277(w_025_277, w_016_001);
  and2 I025_279(w_025_279, w_012_248, w_023_327);
  nand2 I025_282(w_025_282, w_018_019, w_005_000);
  not1 I025_285(w_025_285, w_012_227);
  nand2 I025_287(w_025_287, w_006_000, w_016_019);
  or2  I025_288(w_025_288, w_010_423, w_012_295);
  or2  I025_293(w_025_293, w_002_013, w_023_009);
  nand2 I025_295(w_025_295, w_020_103, w_000_191);
  or2  I025_297(w_025_297, w_007_228, w_018_104);
  and2 I025_311(w_025_311, w_002_010, w_001_003);
  and2 I025_315(w_025_315, w_006_000, w_000_252);
  or2  I025_318(w_025_318, w_023_120, w_010_325);
  and2 I025_320(w_025_320, w_005_208, w_022_103);
  or2  I025_321(w_025_321, w_011_269, w_016_169);
  nand2 I025_322(w_025_322, w_018_098, w_009_172);
  nand2 I025_325(w_025_325, w_013_144, w_014_217);
  and2 I025_326(w_025_326, w_002_007, w_023_034);
  or2  I025_331(w_025_331, w_017_024, w_013_038);
  not1 I025_333(w_025_333, w_019_010);
  or2  I025_336(w_025_336, w_013_239, w_007_032);
  not1 I025_340(w_025_340, w_000_210);
  and2 I025_349(w_025_349, w_006_000, w_022_000);
  and2 I025_350(w_025_350, w_009_234, w_008_106);
  and2 I025_354(w_025_354, w_013_053, w_002_016);
  and2 I025_359(w_025_359, w_014_202, w_023_063);
  and2 I025_362(w_025_362, w_004_465, w_004_405);
  and2 I025_373(w_025_373, w_008_273, w_015_058);
  not1 I025_375(w_025_375, w_003_028);
  and2 I025_376(w_025_376, w_007_003, w_018_123);
  or2  I025_380(w_025_380, w_012_109, w_006_000);
  not1 I025_385(w_025_385, w_009_154);
  and2 I025_388(w_025_388, w_002_014, w_012_007);
  not1 I025_391(w_025_391, w_019_020);
  not1 I025_394(w_025_394, w_008_203);
  nand2 I025_396(w_025_396, w_013_068, w_010_033);
  or2  I025_402(w_025_402, w_009_191, w_017_081);
  nand2 I025_404(w_025_404, w_016_009, w_009_067);
  not1 I025_413(w_025_413, w_007_298);
  and2 I025_416(w_025_416, w_006_000, w_022_145);
  or2  I025_420(w_025_420, w_008_109, w_006_000);
  or2  I025_422(w_025_422, w_013_027, w_015_064);
  nand2 I025_423(w_025_423, w_024_058, w_022_059);
  and2 I025_424(w_025_424, w_011_102, w_001_001);
  not1 I025_428(w_025_428, w_009_137);
  or2  I025_429(w_025_429, w_001_003, w_005_250);
  not1 I025_431(w_025_431, w_004_267);
  nand2 I025_445(w_025_445, w_016_364, w_024_122);
  nand2 I025_446(w_025_446, w_014_185, w_015_069);
  and2 I025_450(w_025_450, w_020_117, w_011_111);
  nand2 I025_456(w_025_456, w_009_136, w_024_197);
  and2 I025_459(w_025_459, w_023_190, w_006_000);
  and2 I025_463(w_025_463, w_005_175, w_008_025);
  nand2 I025_466(w_025_466, w_020_011, w_005_095);
  and2 I025_470(w_025_470, w_014_167, w_023_176);
  not1 I025_471(w_025_471, w_000_262);
  or2  I025_472(w_025_472, w_004_373, w_019_017);
  nand2 I025_476(w_025_476, w_012_108, w_015_028);
  nand2 I025_477(w_025_477, w_006_000, w_017_075);
  not1 I026_002(w_026_002, w_025_070);
  and2 I026_003(w_026_003, w_021_103, w_010_041);
  and2 I026_004(w_026_004, w_016_152, w_013_217);
  nand2 I026_007(w_026_007, w_025_160, w_008_092);
  not1 I026_011(w_026_011, w_007_077);
  or2  I026_012(w_026_012, w_005_121, w_018_078);
  and2 I026_013(w_026_013, w_007_249, w_020_100);
  or2  I026_014(w_026_014, w_003_061, w_004_107);
  or2  I026_017(w_026_017, w_001_001, w_022_057);
  and2 I026_018(w_026_018, w_017_128, w_001_001);
  not1 I026_020(w_026_020, w_007_048);
  or2  I026_021(w_026_021, w_002_020, w_006_000);
  and2 I026_022(w_026_022, w_014_013, w_005_021);
  and2 I026_025(w_026_025, w_011_125, w_020_097);
  not1 I026_033(w_026_033, w_014_016);
  not1 I026_034(w_026_034, w_020_183);
  not1 I026_035(w_026_035, w_008_109);
  not1 I026_036(w_026_036, w_014_240);
  nand2 I026_038(w_026_038, w_007_174, w_011_038);
  not1 I026_039(w_026_039, w_002_007);
  nand2 I026_042(w_026_042, w_011_303, w_021_053);
  nand2 I026_048(w_026_048, w_019_011, w_013_088);
  and2 I026_049(w_026_049, w_008_028, w_020_114);
  not1 I026_050(w_026_050, w_025_155);
  not1 I026_056(w_026_056, w_021_002);
  or2  I026_058(w_026_058, w_018_139, w_006_000);
  and2 I026_060(w_026_060, w_017_177, w_000_400);
  nand2 I026_066(w_026_066, w_015_001, w_018_053);
  nand2 I026_068(w_026_068, w_022_040, w_014_254);
  and2 I026_070(w_026_070, w_023_374, w_023_275);
  and2 I026_072(w_026_072, w_003_036, w_023_110);
  or2  I026_073(w_026_073, w_015_027, w_024_150);
  nand2 I026_082(w_026_082, w_025_069, w_025_373);
  and2 I026_084(w_026_084, w_002_025, w_006_000);
  nand2 I026_087(w_026_087, w_014_081, w_018_132);
  and2 I026_088(w_026_088, w_003_051, w_001_000);
  nand2 I026_091(w_026_091, w_004_215, w_010_404);
  and2 I026_098(w_026_098, w_021_052, w_009_221);
  nand2 I026_099(w_026_099, w_006_000, w_013_180);
  nand2 I026_102(w_026_102, w_017_028, w_005_061);
  not1 I026_103(w_026_103, w_014_014);
  and2 I026_104(w_026_104, w_002_017, w_001_002);
  not1 I026_105(w_026_105, w_022_144);
  or2  I026_113(w_026_113, w_024_004, w_007_317);
  nand2 I026_114(w_026_114, w_000_348, w_011_080);
  and2 I026_118(w_026_118, w_001_004, w_010_357);
  nand2 I026_125(w_026_125, w_007_057, w_023_182);
  nand2 I026_127(w_026_127, w_021_012, w_013_264);
  not1 I026_128(w_026_128, w_009_086);
  or2  I026_131(w_026_131, w_020_125, w_003_037);
  nand2 I026_133(w_026_133, w_014_011, w_025_295);
  and2 I026_137(w_026_137, w_020_126, w_022_084);
  nand2 I026_142(w_026_142, w_009_167, w_020_055);
  not1 I026_145(w_026_145, w_019_034);
  or2  I026_148(w_026_148, w_020_073, w_013_095);
  or2  I026_150(w_026_150, w_008_226, w_000_118);
  or2  I026_151(w_026_151, w_010_176, w_017_109);
  nand2 I026_162(w_026_162, w_019_047, w_005_077);
  not1 I026_173(w_026_173, w_016_375);
  not1 I026_175(w_026_175, w_000_309);
  or2  I026_180(w_026_180, w_024_226, w_003_091);
  nand2 I026_187(w_026_187, w_008_190, w_010_083);
  and2 I026_188(w_026_188, w_009_220, w_014_001);
  nand2 I026_189(w_026_189, w_019_036, w_010_260);
  not1 I026_192(w_026_192, w_010_287);
  not1 I026_193(w_026_193, w_025_402);
  and2 I026_197(w_026_197, w_013_194, w_005_081);
  or2  I026_201(w_026_201, w_006_000, w_009_175);
  or2  I026_204(w_026_204, w_005_022, w_002_012);
  not1 I026_206(w_026_206, w_020_086);
  or2  I026_209(w_026_209, w_006_000, w_014_023);
  or2  I026_210(w_026_210, w_000_348, w_010_175);
  not1 I026_212(w_026_212, w_008_052);
  nand2 I026_213(w_026_213, w_012_004, w_017_092);
  and2 I026_214(w_026_214, w_022_042, w_022_103);
  or2  I026_219(w_026_219, w_019_005, w_002_017);
  and2 I026_227(w_026_227, w_009_168, w_000_280);
  nand2 I026_230(w_026_230, w_017_156, w_006_000);
  nand2 I026_232(w_026_232, w_007_049, w_011_273);
  nand2 I026_242(w_026_242, w_000_445, w_000_171);
  or2  I026_248(w_026_248, w_010_024, w_016_107);
  or2  I026_250(w_026_250, w_007_068, w_002_000);
  not1 I026_251(w_026_251, w_006_000);
  and2 I026_256(w_026_256, w_013_061, w_009_005);
  nand2 I026_260(w_026_260, w_025_471, w_000_101);
  and2 I026_266(w_026_266, w_024_060, w_003_006);
  nand2 I026_268(w_026_268, w_011_318, w_013_066);
  or2  I026_276(w_026_276, w_000_214, w_021_086);
  nand2 I026_280(w_026_280, w_010_316, w_022_056);
  not1 I026_283(w_026_283, w_020_040);
  or2  I026_287(w_026_287, w_005_101, w_012_063);
  not1 I026_294(w_026_294, w_010_425);
  not1 I026_302(w_026_302, w_002_015);
  nand2 I026_305(w_026_305, w_015_043, w_020_016);
  and2 I026_316(w_026_316, w_001_006, w_017_185);
  or2  I026_326(w_026_326, w_024_127, w_014_212);
  or2  I026_328(w_026_328, w_022_071, w_022_148);
  or2  I026_332(w_026_332, w_005_093, w_022_002);
  nand2 I026_334(w_026_334, w_025_466, w_005_228);
  or2  I026_341(w_026_341, w_019_004, w_002_018);
  and2 I026_342(w_026_342, w_012_220, w_016_014);
  nand2 I026_345(w_026_345, w_010_286, w_004_331);
  nand2 I026_346(w_026_346, w_022_007, w_005_011);
  nand2 I026_355(w_026_355, w_024_117, w_016_378);
  nand2 I026_359(w_026_359, w_011_218, w_021_064);
  nand2 I026_361(w_026_361, w_024_090, w_009_086);
  or2  I026_362(w_026_362, w_020_068, w_004_315);
  nand2 I026_363(w_026_363, w_019_013, w_017_081);
  nand2 I026_367(w_026_367, w_010_146, w_024_045);
  not1 I026_370(w_026_370, w_004_202);
  not1 I026_372(w_026_372, w_001_000);
  and2 I026_375(w_026_375, w_007_095, w_017_023);
  and2 I026_377(w_026_377, w_021_048, w_002_024);
  not1 I026_378(w_026_378, w_005_160);
  or2  I026_384(w_026_384, w_011_001, w_024_188);
  or2  I026_386(w_026_386, w_015_078, w_013_046);
  not1 I026_387(w_026_387, w_000_165);
  and2 I026_389(w_026_389, w_020_043, w_025_073);
  nand2 I026_392(w_026_392, w_008_054, w_016_241);
  or2  I027_001(w_027_001, w_019_022, w_005_005);
  or2  I027_004(w_027_004, w_016_248, w_012_040);
  and2 I027_005(w_027_005, w_020_106, w_019_033);
  nand2 I027_006(w_027_006, w_010_382, w_024_057);
  and2 I027_007(w_027_007, w_022_005, w_000_113);
  nand2 I027_008(w_027_008, w_007_390, w_006_000);
  or2  I027_009(w_027_009, w_004_039, w_024_066);
  and2 I027_010(w_027_010, w_003_064, w_003_075);
  or2  I027_011(w_027_011, w_023_028, w_001_003);
  nand2 I027_014(w_027_014, w_007_255, w_004_038);
  nand2 I027_018(w_027_018, w_010_131, w_000_233);
  and2 I027_019(w_027_019, w_013_087, w_018_012);
  not1 I027_020(w_027_020, w_014_170);
  and2 I027_022(w_027_022, w_002_025, w_026_070);
  and2 I027_025(w_027_025, w_021_032, w_020_108);
  and2 I027_027(w_027_027, w_003_066, w_012_040);
  not1 I027_028(w_027_028, w_005_094);
  nand2 I027_030(w_027_030, w_005_203, w_001_004);
  not1 I027_031(w_027_031, w_014_005);
  nand2 I027_032(w_027_032, w_020_024, w_006_000);
  and2 I027_033(w_027_033, w_009_113, w_024_124);
  not1 I027_035(w_027_035, w_012_161);
  and2 I027_039(w_027_039, w_014_159, w_003_067);
  or2  I027_041(w_027_041, w_004_183, w_020_012);
  nand2 I027_042(w_027_042, w_014_231, w_014_014);
  nand2 I027_057(w_027_057, w_002_000, w_011_069);
  and2 I027_060(w_027_060, w_001_000, w_002_008);
  nand2 I027_063(w_027_063, w_010_318, w_022_079);
  not1 I027_064(w_027_064, w_006_000);
  and2 I027_067(w_027_067, w_016_197, w_018_160);
  not1 I027_069(w_027_069, w_003_100);
  nand2 I027_070(w_027_070, w_023_307, w_013_089);
  not1 I027_074(w_027_074, w_014_005);
  nand2 I027_075(w_027_075, w_020_060, w_017_053);
  or2  I027_076(w_027_076, w_020_153, w_006_000);
  and2 I027_080(w_027_080, w_022_084, w_010_049);
  not1 I027_086(w_027_086, w_009_125);
  and2 I027_088(w_027_088, w_000_447, w_018_074);
  or2  I027_091(w_027_091, w_010_044, w_009_035);
  or2  I027_101(w_027_101, w_016_178, w_018_015);
  or2  I027_104(w_027_104, w_012_138, w_020_078);
  not1 I027_108(w_027_108, w_026_188);
  nand2 I027_111(w_027_111, w_007_390, w_001_005);
  or2  I027_112(w_027_112, w_014_165, w_019_000);
  or2  I027_114(w_027_114, w_013_101, w_017_030);
  or2  I027_115(w_027_115, w_017_027, w_022_107);
  not1 I027_120(w_027_120, w_009_159);
  or2  I027_123(w_027_123, w_009_170, w_020_150);
  not1 I027_128(w_027_128, w_005_228);
  and2 I027_133(w_027_133, w_005_221, w_000_377);
  nand2 I027_134(w_027_134, w_008_092, w_008_225);
  nand2 I027_135(w_027_135, w_003_043, w_020_079);
  not1 I027_138(w_027_138, w_017_020);
  and2 I027_141(w_027_141, w_020_034, w_017_083);
  and2 I027_147(w_027_147, w_018_047, w_013_223);
  or2  I027_150(w_027_150, w_008_023, w_021_108);
  or2  I027_152(w_027_152, w_004_292, w_006_000);
  not1 I027_153(w_027_153, w_023_314);
  or2  I027_154(w_027_154, w_010_037, w_003_081);
  nand2 I027_155(w_027_155, w_010_079, w_002_012);
  nand2 I027_163(w_027_163, w_021_014, w_006_000);
  nand2 I027_165(w_027_165, w_017_099, w_004_320);
  and2 I027_166(w_027_166, w_022_141, w_014_125);
  and2 I027_168(w_027_168, w_025_194, w_001_006);
  nand2 I027_169(w_027_169, w_001_000, w_014_161);
  and2 I027_172(w_027_172, w_026_392, w_013_018);
  and2 I027_175(w_027_175, w_004_240, w_000_250);
  not1 I027_178(w_027_178, w_017_060);
  and2 I027_183(w_027_183, w_015_105, w_002_003);
  and2 I027_184(w_027_184, w_005_171, w_003_068);
  not1 I027_185(w_027_185, w_009_024);
  or2  I027_186(w_027_186, w_025_020, w_022_062);
  or2  I027_194(w_027_194, w_010_196, w_001_002);
  or2  I027_196(w_027_196, w_014_092, w_017_063);
  nand2 I027_198(w_027_198, w_021_049, w_001_003);
  not1 I027_199(w_027_199, w_024_277);
  and2 I027_201(w_027_201, w_018_083, w_008_127);
  and2 I027_203(w_027_203, w_004_283, w_021_027);
  not1 I027_209(w_027_209, w_016_287);
  or2  I027_211(w_027_211, w_022_156, w_015_036);
  nand2 I027_215(w_027_215, w_010_327, w_024_078);
  nand2 I027_217(w_027_217, w_024_280, w_022_069);
  or2  I027_218(w_027_218, w_006_000, w_008_066);
  not1 I027_226(w_027_226, w_009_030);
  and2 I027_228(w_027_228, w_014_141, w_013_185);
  nand2 I027_232(w_027_232, w_016_384, w_019_010);
  and2 I027_235(w_027_235, w_007_309, w_011_067);
  not1 I027_237(w_027_237, w_023_401);
  and2 I027_239(w_027_239, w_008_153, w_024_151);
  nand2 I027_240(w_027_240, w_005_214, w_020_013);
  and2 I027_241(w_027_241, w_023_400, w_013_133);
  or2  I027_242(w_027_242, w_020_069, w_008_005);
  nand2 I027_249(w_027_249, w_009_224, w_005_017);
  nand2 I027_251(w_027_251, w_025_066, w_017_117);
  and2 I027_256(w_027_256, w_010_262, w_016_369);
  or2  I027_257(w_027_257, w_022_011, w_005_195);
  and2 I027_258(w_027_258, w_022_005, w_008_103);
  not1 I027_262(w_027_262, w_010_384);
  nand2 I027_263(w_027_263, w_020_124, w_015_090);
  nand2 I027_264(w_027_264, w_011_063, w_008_202);
  and2 I027_268(w_027_268, w_024_189, w_003_084);
  or2  I027_275(w_027_275, w_010_291, w_002_025);
  not1 I027_278(w_027_278, w_007_136);
  not1 I027_280(w_027_280, w_003_046);
  and2 I027_282(w_027_282, w_024_090, w_009_052);
  and2 I027_287(w_027_287, w_019_048, w_003_050);
  and2 I027_295(w_027_295, w_006_000, w_022_079);
  and2 I027_299(w_027_299, w_002_021, w_014_161);
  nand2 I027_312(w_027_312, w_012_325, w_004_290);
  nand2 I027_313(w_027_313, w_003_062, w_000_350);
  not1 I027_321(w_027_321, w_001_003);
  or2  I027_324(w_027_324, w_014_053, w_014_209);
  and2 I027_325(w_027_325, w_008_244, w_018_026);
  nand2 I027_328(w_027_328, w_001_002, w_019_010);
  or2  I027_329(w_027_329, w_019_038, w_005_119);
  nand2 I027_331(w_027_331, w_009_140, w_013_191);
  not1 I027_332(w_027_332, w_004_385);
  or2  I027_337(w_027_337, w_011_019, w_001_000);
  not1 I027_339(w_027_339, w_010_151);
  nand2 I027_341(w_027_341, w_002_005, w_006_000);
  not1 I027_347(w_027_347, w_017_176);
  or2  I027_348(w_027_348, w_020_013, w_018_071);
  not1 I027_354(w_027_354, w_005_142);
  nand2 I027_355(w_027_355, w_025_095, w_025_459);
  nand2 I027_357(w_027_357, w_009_091, w_007_305);
  not1 I027_359(w_027_359, w_020_156);
  not1 I027_362(w_027_362, w_008_004);
  and2 I027_366(w_027_366, w_014_092, w_005_101);
  or2  I027_367(w_027_367, w_023_185, w_015_026);
  or2  I027_370(w_027_370, w_009_003, w_013_036);
  not1 I027_372(w_027_372, w_007_027);
  and2 I027_378(w_027_378, w_009_176, w_020_074);
  nand2 I027_382(w_027_382, w_008_093, w_025_082);
  nand2 I027_389(w_027_389, w_010_344, w_001_001);
  nand2 I027_394(w_027_394, w_018_039, w_011_291);
  and2 I027_400(w_027_400, w_011_039, w_023_059);
  or2  I027_403(w_027_403, w_013_066, w_011_333);
  not1 I027_404(w_027_404, w_011_043);
  not1 I027_412(w_027_412, w_024_067);
  nand2 I027_416(w_027_416, w_013_166, w_000_195);
  and2 I027_426(w_027_426, w_007_271, w_013_093);
  and2 I027_427(w_027_427, w_000_411, w_023_104);
  nand2 I027_431(w_027_431, w_007_268, w_003_046);
  and2 I027_438(w_027_438, w_022_158, w_018_006);
  or2  I027_439(w_027_439, w_019_000, w_013_043);
  not1 I027_443(w_027_443, w_018_100);
  nand2 I027_444(w_027_444, w_015_090, w_025_150);
  nand2 I027_449(w_027_449, w_005_176, w_015_073);
  nand2 I027_452(w_027_452, w_006_000, w_012_144);
  nand2 I028_000(w_028_000, w_010_201, w_024_241);
  or2  I028_001(w_028_001, w_001_002, w_027_426);
  and2 I028_004(w_028_004, w_018_002, w_019_007);
  and2 I028_005(w_028_005, w_005_070, w_024_136);
  and2 I028_006(w_028_006, w_017_020, w_003_031);
  or2  I028_008(w_028_008, w_005_154, w_027_237);
  not1 I028_009(w_028_009, w_008_198);
  and2 I028_011(w_028_011, w_007_261, w_012_368);
  and2 I028_013(w_028_013, w_012_189, w_025_340);
  or2  I028_014(w_028_014, w_004_321, w_006_000);
  and2 I028_015(w_028_015, w_006_000, w_009_022);
  nand2 I028_016(w_028_016, w_020_146, w_023_324);
  and2 I028_017(w_028_017, w_016_372, w_017_116);
  and2 I028_019(w_028_019, w_000_399, w_024_033);
  nand2 I028_029(w_028_029, w_006_000, w_019_023);
  or2  I028_032(w_028_032, w_001_005, w_002_014);
  not1 I028_035(w_028_035, w_025_385);
  and2 I028_039(w_028_039, w_005_057, w_002_023);
  or2  I028_040(w_028_040, w_000_232, w_014_197);
  or2  I028_041(w_028_041, w_023_163, w_023_063);
  not1 I028_042(w_028_042, w_004_363);
  nand2 I028_047(w_028_047, w_016_027, w_012_379);
  not1 I028_048(w_028_048, w_007_210);
  and2 I028_049(w_028_049, w_011_082, w_001_003);
  nand2 I028_052(w_028_052, w_009_118, w_024_032);
  or2  I028_056(w_028_056, w_022_102, w_024_132);
  or2  I028_058(w_028_058, w_010_368, w_020_120);
  not1 I028_060(w_028_060, w_009_016);
  not1 I028_070(w_028_070, w_017_014);
  and2 I028_073(w_028_073, w_010_041, w_024_229);
  nand2 I028_074(w_028_074, w_016_099, w_014_131);
  or2  I028_076(w_028_076, w_007_156, w_003_086);
  or2  I028_082(w_028_082, w_004_318, w_006_000);
  not1 I028_083(w_028_083, w_009_229);
  or2  I028_084(w_028_084, w_025_394, w_022_138);
  nand2 I028_085(w_028_085, w_008_175, w_023_059);
  nand2 I028_087(w_028_087, w_019_021, w_020_145);
  nand2 I028_096(w_028_096, w_010_134, w_009_033);
  not1 I028_100(w_028_100, w_004_371);
  not1 I028_108(w_028_108, w_011_301);
  nand2 I028_109(w_028_109, w_020_112, w_019_010);
  and2 I028_115(w_028_115, w_010_273, w_027_275);
  and2 I028_118(w_028_118, w_002_024, w_017_081);
  not1 I028_119(w_028_119, w_000_389);
  not1 I028_123(w_028_123, w_010_172);
  nand2 I028_128(w_028_128, w_014_125, w_016_091);
  and2 I028_129(w_028_129, w_024_018, w_003_072);
  or2  I028_130(w_028_130, w_013_152, w_011_192);
  not1 I028_132(w_028_132, w_015_085);
  not1 I028_144(w_028_144, w_001_003);
  not1 I028_149(w_028_149, w_009_063);
  or2  I028_151(w_028_151, w_020_032, w_014_222);
  and2 I028_159(w_028_159, w_015_082, w_012_303);
  and2 I028_171(w_028_171, w_025_091, w_027_295);
  and2 I028_174(w_028_174, w_015_129, w_006_000);
  nand2 I028_184(w_028_184, w_001_000, w_024_240);
  and2 I028_187(w_028_187, w_024_169, w_011_124);
  not1 I028_188(w_028_188, w_027_280);
  or2  I028_197(w_028_197, w_024_059, w_019_001);
  and2 I028_199(w_028_199, w_001_001, w_012_353);
  or2  I028_200(w_028_200, w_002_015, w_024_112);
  not1 I028_201(w_028_201, w_023_256);
  and2 I028_205(w_028_205, w_026_060, w_013_246);
  or2  I028_206(w_028_206, w_019_022, w_001_002);
  or2  I028_208(w_028_208, w_023_330, w_019_012);
  not1 I028_215(w_028_215, w_023_018);
  not1 I028_216(w_028_216, w_009_146);
  and2 I028_221(w_028_221, w_007_004, w_006_000);
  not1 I028_232(w_028_232, w_023_220);
  nand2 I028_236(w_028_236, w_016_076, w_026_250);
  or2  I028_237(w_028_237, w_016_280, w_006_000);
  and2 I028_239(w_028_239, w_008_001, w_017_020);
  not1 I028_241(w_028_241, w_006_000);
  not1 I028_254(w_028_254, w_024_065);
  not1 I028_255(w_028_255, w_026_173);
  nand2 I028_258(w_028_258, w_023_309, w_009_107);
  and2 I028_262(w_028_262, w_021_023, w_013_040);
  or2  I028_266(w_028_266, w_004_243, w_004_156);
  nand2 I028_267(w_028_267, w_003_017, w_025_394);
  nand2 I028_268(w_028_268, w_017_135, w_018_168);
  and2 I028_270(w_028_270, w_011_016, w_003_077);
  and2 I028_277(w_028_277, w_007_016, w_023_196);
  not1 I028_284(w_028_284, w_003_043);
  and2 I028_290(w_028_290, w_006_000, w_014_163);
  or2  I028_292(w_028_292, w_020_000, w_013_068);
  not1 I028_296(w_028_296, w_019_035);
  or2  I028_299(w_028_299, w_019_035, w_006_000);
  not1 I028_305(w_028_305, w_020_049);
  nand2 I028_308(w_028_308, w_006_000, w_026_020);
  and2 I028_309(w_028_309, w_024_170, w_002_019);
  nand2 I028_313(w_028_313, w_012_055, w_005_021);
  or2  I028_316(w_028_316, w_008_004, w_006_000);
  and2 I028_323(w_028_323, w_008_152, w_022_006);
  or2  I028_324(w_028_324, w_001_002, w_011_309);
  and2 I028_325(w_028_325, w_008_082, w_010_288);
  and2 I028_332(w_028_332, w_011_144, w_000_450);
  not1 I028_334(w_028_334, w_016_164);
  or2  I028_335(w_028_335, w_018_017, w_014_196);
  nand2 I028_339(w_028_339, w_005_173, w_012_255);
  and2 I028_341(w_028_341, w_008_017, w_004_102);
  nand2 I028_345(w_028_345, w_006_000, w_025_391);
  not1 I028_348(w_028_348, w_004_194);
  nand2 I028_350(w_028_350, w_012_004, w_013_193);
  nand2 I028_353(w_028_353, w_022_117, w_002_005);
  or2  I028_355(w_028_355, w_013_039, w_015_124);
  nand2 I028_356(w_028_356, w_027_264, w_011_089);
  or2  I028_360(w_028_360, w_016_371, w_016_214);
  or2  I028_364(w_028_364, w_001_005, w_025_074);
  not1 I028_370(w_028_370, w_017_026);
  not1 I028_379(w_028_379, w_007_147);
  not1 I028_381(w_028_381, w_014_116);
  and2 I028_382(w_028_382, w_020_015, w_023_306);
  not1 I028_386(w_028_386, w_000_385);
  or2  I028_395(w_028_395, w_010_400, w_003_085);
  and2 I028_397(w_028_397, w_003_064, w_025_315);
  and2 I029_001(w_029_001, w_007_193, w_008_191);
  and2 I029_006(w_029_006, w_014_013, w_007_366);
  or2  I029_010(w_029_010, w_018_124, w_027_030);
  or2  I029_012(w_029_012, w_015_007, w_021_089);
  or2  I029_013(w_029_013, w_021_048, w_016_345);
  and2 I029_014(w_029_014, w_028_073, w_027_152);
  or2  I029_017(w_029_017, w_009_043, w_026_384);
  or2  I029_019(w_029_019, w_023_267, w_015_002);
  nand2 I029_024(w_029_024, w_001_000, w_017_101);
  or2  I029_025(w_029_025, w_019_045, w_011_312);
  or2  I029_028(w_029_028, w_004_301, w_015_074);
  not1 I029_029(w_029_029, w_019_014);
  or2  I029_031(w_029_031, w_024_054, w_020_182);
  not1 I029_039(w_029_039, w_014_009);
  nand2 I029_040(w_029_040, w_016_068, w_018_124);
  nand2 I029_043(w_029_043, w_018_160, w_017_077);
  not1 I029_044(w_029_044, w_027_431);
  not1 I029_045(w_029_045, w_006_000);
  and2 I029_047(w_029_047, w_008_077, w_018_163);
  or2  I029_052(w_029_052, w_002_024, w_020_115);
  or2  I029_057(w_029_057, w_004_005, w_013_124);
  and2 I029_059(w_029_059, w_026_378, w_018_243);
  nand2 I029_061(w_029_061, w_005_001, w_017_058);
  or2  I029_063(w_029_063, w_014_008, w_020_154);
  nand2 I029_067(w_029_067, w_016_191, w_019_011);
  not1 I029_068(w_029_068, w_025_260);
  nand2 I029_071(w_029_071, w_018_186, w_018_142);
  nand2 I029_073(w_029_073, w_016_257, w_015_082);
  nand2 I029_075(w_029_075, w_019_019, w_025_245);
  and2 I029_077(w_029_077, w_024_116, w_014_131);
  nand2 I029_078(w_029_078, w_013_232, w_026_003);
  nand2 I029_080(w_029_080, w_001_006, w_014_161);
  and2 I029_082(w_029_082, w_003_072, w_006_000);
  and2 I029_083(w_029_083, w_016_153, w_000_451);
  or2  I029_086(w_029_086, w_026_099, w_007_006);
  and2 I029_095(w_029_095, w_005_144, w_002_015);
  or2  I029_096(w_029_096, w_000_370, w_028_200);
  or2  I029_097(w_029_097, w_012_063, w_004_186);
  not1 I029_098(w_029_098, w_010_004);
  and2 I029_099(w_029_099, w_026_287, w_025_326);
  and2 I029_107(w_029_107, w_016_374, w_026_268);
  or2  I029_111(w_029_111, w_028_355, w_025_149);
  not1 I029_112(w_029_112, w_007_266);
  or2  I029_113(w_029_113, w_023_209, w_024_266);
  or2  I029_115(w_029_115, w_005_196, w_008_008);
  nand2 I029_116(w_029_116, w_016_233, w_016_223);
  not1 I029_118(w_029_118, w_013_146);
  and2 I029_119(w_029_119, w_002_014, w_010_151);
  nand2 I029_121(w_029_121, w_002_021, w_006_000);
  not1 I029_122(w_029_122, w_006_000);
  and2 I029_124(w_029_124, w_020_091, w_002_014);
  not1 I029_128(w_029_128, w_001_002);
  not1 I029_130(w_029_130, w_019_011);
  not1 I029_133(w_029_133, w_005_236);
  and2 I029_136(w_029_136, w_007_124, w_020_043);
  or2  I029_137(w_029_137, w_013_007, w_007_046);
  not1 I029_139(w_029_139, w_028_316);
  or2  I029_141(w_029_141, w_006_000, w_021_018);
  and2 I029_142(w_029_142, w_025_106, w_028_397);
  nand2 I029_147(w_029_147, w_009_084, w_018_020);
  and2 I029_149(w_029_149, w_002_027, w_027_175);
  and2 I029_151(w_029_151, w_001_000, w_026_033);
  and2 I029_152(w_029_152, w_024_287, w_007_340);
  nand2 I029_153(w_029_153, w_000_026, w_010_020);
  or2  I029_154(w_029_154, w_010_450, w_005_089);
  and2 I029_157(w_029_157, w_006_000, w_022_142);
  or2  I029_160(w_029_160, w_008_000, w_027_033);
  and2 I029_161(w_029_161, w_015_116, w_013_068);
  nand2 I029_163(w_029_163, w_009_221, w_025_085);
  not1 I029_166(w_029_166, w_027_076);
  or2  I029_167(w_029_167, w_025_063, w_009_059);
  and2 I029_172(w_029_172, w_015_066, w_008_061);
  or2  I029_173(w_029_173, w_006_000, w_017_009);
  and2 I029_175(w_029_175, w_011_071, w_010_121);
  and2 I029_176(w_029_176, w_007_286, w_013_044);
  and2 I029_177(w_029_177, w_025_020, w_023_335);
  not1 I029_178(w_029_178, w_024_078);
  or2  I029_179(w_029_179, w_024_191, w_005_161);
  not1 I029_181(w_029_181, w_002_005);
  not1 I029_182(w_029_182, w_005_087);
  nand2 I029_184(w_029_184, w_007_398, w_013_227);
  not1 I029_186(w_029_186, w_019_036);
  and2 I029_187(w_029_187, w_013_100, w_007_105);
  nand2 I029_188(w_029_188, w_018_068, w_022_041);
  not1 I029_189(w_029_189, w_028_128);
  nand2 I029_192(w_029_192, w_013_189, w_022_013);
  not1 I029_194(w_029_194, w_010_196);
  not1 I029_195(w_029_195, w_024_076);
  not1 I029_197(w_029_197, w_014_091);
  and2 I029_198(w_029_198, w_005_220, w_014_002);
  or2  I029_201(w_029_201, w_015_089, w_018_110);
  nand2 I029_202(w_029_202, w_006_000, w_003_033);
  and2 I029_204(w_029_204, w_001_001, w_011_012);
  or2  I029_213(w_029_213, w_003_090, w_015_022);
  or2  I029_215(w_029_215, w_012_339, w_002_002);
  or2  I029_217(w_029_217, w_009_190, w_001_002);
  and2 I029_220(w_029_220, w_006_000, w_014_009);
  nand2 I029_221(w_029_221, w_022_050, w_015_017);
  nand2 I029_222(w_029_222, w_003_017, w_011_206);
  nand2 I029_223(w_029_223, w_003_019, w_008_162);
  nand2 I029_225(w_029_225, w_001_003, w_027_226);
  or2  I029_229(w_029_229, w_023_013, w_023_290);
  not1 I029_231(w_029_231, w_006_000);
  not1 I029_232(w_029_232, w_024_070);
  and2 I029_233(w_029_233, w_012_165, w_014_027);
  nand2 I029_234(w_029_234, w_022_143, w_028_074);
  nand2 I029_237(w_029_237, w_013_066, w_025_476);
  nand2 I029_240(w_029_240, w_002_007, w_028_323);
  not1 I029_241(w_029_241, w_027_147);
  nand2 I029_242(w_029_242, w_019_010, w_021_079);
  not1 I029_243(w_029_243, w_024_245);
  nand2 I029_245(w_029_245, w_023_052, w_004_199);
  nand2 I029_246(w_029_246, w_021_017, w_021_079);
  and2 I029_247(w_029_247, w_016_230, w_028_267);
  nand2 I029_248(w_029_250, w_008_083, w_029_249);
  not1 I029_249(w_029_251, w_029_250);
  and2 I029_250(w_029_252, w_029_251, w_019_048);
  and2 I029_251(w_029_253, w_029_252, w_012_122);
  not1 I029_252(w_029_254, w_029_253);
  not1 I029_253(w_029_255, w_029_254);
  and2 I029_254(w_029_256, w_029_255, w_029_265);
  or2  I029_255(w_029_249, w_018_000, w_029_256);
  or2  I029_256(w_029_261, w_003_069, w_029_260);
  or2  I029_257(w_029_262, w_028_085, w_029_261);
  or2  I029_258(w_029_263, w_022_131, w_029_262);
  not1 I029_259(w_029_260, w_029_256);
  and2 I029_260(w_029_265, w_020_055, w_029_263);
  not1 I030_002(w_030_002, w_028_119);
  or2  I030_003(w_030_003, w_009_036, w_020_049);
  not1 I030_006(w_030_006, w_003_028);
  or2  I030_010(w_030_010, w_005_106, w_020_137);
  and2 I030_012(w_030_012, w_025_095, w_005_170);
  or2  I030_016(w_030_016, w_020_095, w_018_054);
  not1 I030_017(w_030_017, w_008_020);
  nand2 I030_019(w_030_019, w_009_044, w_024_181);
  nand2 I030_022(w_030_022, w_018_239, w_008_118);
  or2  I030_024(w_030_024, w_026_214, w_008_068);
  and2 I030_026(w_030_026, w_027_416, w_025_276);
  and2 I030_027(w_030_027, w_016_297, w_029_233);
  not1 I030_029(w_030_029, w_021_016);
  not1 I030_030(w_030_030, w_000_279);
  or2  I030_031(w_030_031, w_018_124, w_027_382);
  not1 I030_035(w_030_035, w_018_097);
  and2 I030_040(w_030_040, w_018_014, w_012_201);
  nand2 I030_041(w_030_041, w_012_089, w_005_132);
  not1 I030_043(w_030_043, w_010_332);
  nand2 I030_045(w_030_045, w_009_231, w_013_051);
  and2 I030_047(w_030_047, w_019_047, w_015_115);
  and2 I030_049(w_030_049, w_016_222, w_018_288);
  not1 I030_051(w_030_051, w_026_346);
  or2  I030_053(w_030_053, w_010_427, w_027_069);
  not1 I030_054(w_030_054, w_005_173);
  not1 I030_055(w_030_055, w_018_086);
  nand2 I030_056(w_030_056, w_016_049, w_017_039);
  not1 I030_059(w_030_059, w_019_011);
  nand2 I030_060(w_030_060, w_028_267, w_024_048);
  or2  I030_061(w_030_061, w_023_319, w_017_045);
  and2 I030_062(w_030_062, w_010_108, w_022_075);
  not1 I030_065(w_030_065, w_013_019);
  or2  I030_066(w_030_066, w_025_354, w_018_300);
  not1 I030_067(w_030_067, w_017_035);
  not1 I030_068(w_030_068, w_018_169);
  or2  I030_071(w_030_071, w_012_005, w_001_003);
  nand2 I030_072(w_030_072, w_024_016, w_017_040);
  nand2 I030_076(w_030_076, w_000_338, w_016_058);
  or2  I030_077(w_030_077, w_000_038, w_015_061);
  nand2 I030_078(w_030_078, w_019_005, w_020_125);
  and2 I030_080(w_030_080, w_013_145, w_023_306);
  or2  I030_081(w_030_081, w_015_064, w_025_288);
  and2 I030_085(w_030_085, w_015_044, w_023_121);
  and2 I030_086(w_030_086, w_009_064, w_006_000);
  not1 I030_087(w_030_087, w_013_030);
  not1 I030_088(w_030_088, w_008_318);
  not1 I030_089(w_030_089, w_003_028);
  and2 I030_090(w_030_090, w_022_133, w_016_045);
  not1 I030_091(w_030_091, w_004_025);
  not1 I030_093(w_030_093, w_016_278);
  and2 I030_096(w_030_096, w_004_378, w_024_019);
  nand2 I030_097(w_030_097, w_022_057, w_015_102);
  nand2 I030_098(w_030_098, w_010_192, w_004_256);
  nand2 I030_099(w_030_099, w_008_199, w_016_029);
  or2  I030_101(w_030_101, w_011_087, w_015_020);
  and2 I030_107(w_030_107, w_013_177, w_009_175);
  and2 I030_113(w_030_113, w_020_173, w_020_048);
  not1 I030_116(w_030_116, w_016_263);
  and2 I030_118(w_030_118, w_000_275, w_021_008);
  nand2 I030_119(w_030_119, w_007_298, w_006_000);
  and2 I030_122(w_030_122, w_014_198, w_018_018);
  or2  I030_124(w_030_124, w_021_050, w_015_120);
  and2 I030_128(w_030_128, w_011_186, w_018_256);
  not1 I030_129(w_030_129, w_007_097);
  and2 I030_132(w_030_132, w_006_000, w_029_133);
  nand2 I030_133(w_030_133, w_018_108, w_002_011);
  not1 I030_135(w_030_135, w_025_424);
  or2  I030_136(w_030_136, w_024_072, w_016_394);
  nand2 I030_137(w_030_137, w_003_001, w_010_142);
  or2  I030_138(w_030_138, w_018_075, w_020_054);
  and2 I030_139(w_030_139, w_019_040, w_005_034);
  nand2 I030_140(w_030_140, w_007_319, w_003_012);
  and2 I030_144(w_030_144, w_018_218, w_013_009);
  and2 I030_146(w_030_146, w_009_098, w_007_303);
  not1 I030_147(w_030_147, w_012_143);
  nand2 I030_148(w_030_148, w_020_046, w_021_010);
  not1 I030_150(w_030_150, w_021_078);
  not1 I030_151(w_030_151, w_001_001);
  and2 I030_157(w_030_157, w_017_168, w_005_113);
  nand2 I030_160(w_030_160, w_023_041, w_005_026);
  not1 I030_170(w_030_170, w_012_279);
  or2  I030_172(w_030_172, w_017_122, w_021_027);
  not1 I030_175(w_030_175, w_010_263);
  or2  I030_176(w_030_176, w_015_080, w_020_089);
  or2  I030_178(w_030_178, w_011_214, w_028_290);
  and2 I030_180(w_030_180, w_020_062, w_022_013);
  not1 I030_184(w_030_184, w_027_359);
  nand2 I030_185(w_030_185, w_000_073, w_026_341);
  or2  I030_186(w_030_186, w_007_123, w_016_225);
  or2  I030_188(w_030_188, w_005_156, w_019_022);
  and2 I030_189(w_030_189, w_004_016, w_015_031);
  and2 I030_191(w_030_191, w_021_030, w_027_104);
  and2 I030_193(w_030_193, w_015_120, w_013_194);
  and2 I030_196(w_030_196, w_003_074, w_004_157);
  and2 I030_199(w_030_199, w_001_002, w_012_025);
  nand2 I031_000(w_031_000, w_020_088, w_006_000);
  nand2 I031_001(w_031_001, w_029_187, w_029_246);
  nand2 I031_002(w_031_002, w_027_025, w_015_114);
  or2  I031_003(w_031_003, w_029_136, w_023_039);
  or2  I031_004(w_031_004, w_030_006, w_025_089);
  not1 I031_005(w_031_005, w_015_064);
  not1 I031_006(w_031_006, w_005_098);
  or2  I031_007(w_031_007, w_025_165, w_002_012);
  and2 I031_008(w_031_008, w_030_139, w_024_040);
  or2  I031_010(w_031_010, w_002_025, w_008_056);
  or2  I031_011(w_031_011, w_023_006, w_018_051);
  not1 I031_012(w_031_012, w_022_044);
  and2 I031_013(w_031_013, w_019_016, w_005_154);
  nand2 I031_014(w_031_014, w_028_073, w_007_091);
  or2  I031_015(w_031_015, w_006_000, w_019_038);
  not1 I031_016(w_031_016, w_006_000);
  nand2 I031_017(w_031_017, w_007_283, w_015_015);
  and2 I031_018(w_031_018, w_005_035, w_016_034);
  not1 I031_019(w_031_019, w_005_229);
  not1 I031_020(w_031_020, w_023_228);
  and2 I031_021(w_031_021, w_007_094, w_025_156);
  nand2 I031_022(w_031_022, w_024_294, w_021_027);
  and2 I031_023(w_031_023, w_019_009, w_028_262);
  and2 I031_024(w_031_024, w_004_397, w_015_018);
  or2  I031_025(w_031_025, w_018_306, w_026_050);
  and2 I031_027(w_031_027, w_002_007, w_014_085);
  and2 I031_029(w_031_029, w_001_001, w_006_000);
  not1 I031_030(w_031_030, w_004_445);
  nand2 I031_031(w_031_031, w_017_123, w_003_009);
  or2  I031_032(w_031_032, w_029_115, w_009_038);
  nand2 I031_033(w_031_033, w_010_135, w_016_385);
  not1 I031_034(w_031_034, w_030_122);
  nand2 I031_036(w_031_036, w_017_067, w_001_001);
  and2 I031_037(w_031_037, w_028_083, w_013_152);
  and2 I031_038(w_031_038, w_030_067, w_027_163);
  or2  I031_040(w_031_040, w_024_025, w_006_000);
  nand2 I031_041(w_031_041, w_006_000, w_018_105);
  nand2 I031_042(w_031_042, w_019_012, w_006_000);
  or2  I031_043(w_031_043, w_013_205, w_011_333);
  not1 I031_044(w_031_044, w_003_079);
  not1 I031_045(w_031_045, w_028_299);
  not1 I031_046(w_031_046, w_021_077);
  nand2 I031_048(w_031_048, w_005_238, w_003_096);
  and2 I031_049(w_031_049, w_004_433, w_018_153);
  and2 I031_050(w_031_050, w_006_000, w_027_014);
  and2 I031_051(w_031_051, w_023_140, w_011_128);
  not1 I031_052(w_031_052, w_008_081);
  or2  I031_053(w_031_053, w_027_357, w_027_010);
  and2 I031_054(w_031_054, w_028_397, w_000_452);
  and2 I031_055(w_031_055, w_002_017, w_008_103);
  nand2 I031_056(w_031_056, w_026_102, w_003_020);
  or2  I031_057(w_031_057, w_030_136, w_002_020);
  or2  I031_058(w_031_058, w_013_253, w_010_347);
  not1 I031_061(w_031_061, w_024_075);
  and2 I031_062(w_031_062, w_001_003, w_017_046);
  not1 I031_063(w_031_063, w_018_212);
  nand2 I031_064(w_031_064, w_018_026, w_009_140);
  not1 I031_065(w_031_065, w_022_131);
  or2  I031_066(w_031_066, w_009_164, w_008_125);
  or2  I031_067(w_031_067, w_000_179, w_018_107);
  and2 I032_000(w_032_000, w_013_011, w_003_097);
  not1 I032_002(w_032_002, w_014_225);
  and2 I032_003(w_032_003, w_015_046, w_023_269);
  nand2 I032_004(w_032_004, w_022_018, w_012_114);
  nand2 I032_006(w_032_006, w_030_024, w_019_047);
  and2 I032_008(w_032_008, w_013_006, w_027_111);
  nand2 I032_011(w_032_011, w_026_068, w_023_350);
  not1 I032_013(w_032_013, w_029_044);
  not1 I032_014(w_032_014, w_019_040);
  not1 I032_015(w_032_015, w_008_131);
  or2  I032_018(w_032_018, w_023_180, w_030_170);
  not1 I032_019(w_032_019, w_014_070);
  or2  I032_022(w_032_022, w_013_167, w_010_041);
  not1 I032_023(w_032_023, w_009_174);
  and2 I032_025(w_032_025, w_027_064, w_003_012);
  not1 I032_026(w_032_026, w_017_154);
  and2 I032_027(w_032_027, w_023_239, w_021_108);
  nand2 I032_030(w_032_030, w_010_107, w_016_310);
  or2  I032_034(w_032_034, w_002_013, w_001_006);
  nand2 I032_035(w_032_035, w_030_191, w_027_209);
  or2  I032_037(w_032_037, w_016_073, w_003_044);
  and2 I032_039(w_032_039, w_025_180, w_001_006);
  not1 I032_041(w_032_041, w_014_234);
  or2  I032_042(w_032_042, w_012_125, w_024_072);
  not1 I032_043(w_032_043, w_021_031);
  not1 I032_045(w_032_045, w_009_232);
  and2 I032_048(w_032_048, w_022_117, w_013_150);
  nand2 I032_049(w_032_049, w_007_109, w_005_228);
  not1 I032_051(w_032_051, w_030_030);
  not1 I032_052(w_032_052, w_031_064);
  nand2 I032_053(w_032_053, w_003_049, w_006_000);
  not1 I032_054(w_032_054, w_014_193);
  or2  I032_055(w_032_055, w_023_354, w_020_182);
  or2  I032_058(w_032_058, w_019_016, w_021_025);
  nand2 I032_059(w_032_059, w_024_295, w_022_116);
  or2  I032_061(w_032_061, w_030_133, w_031_031);
  and2 I032_065(w_032_065, w_012_138, w_031_020);
  or2  I032_066(w_032_066, w_021_000, w_004_395);
  or2  I032_068(w_032_068, w_028_001, w_002_027);
  or2  I032_069(w_032_069, w_007_209, w_012_046);
  nand2 I032_070(w_032_070, w_001_004, w_003_050);
  nand2 I032_071(w_032_071, w_011_300, w_017_114);
  and2 I032_072(w_032_072, w_010_359, w_004_142);
  nand2 I032_073(w_032_073, w_016_095, w_028_262);
  and2 I032_074(w_032_074, w_005_125, w_003_036);
  nand2 I032_077(w_032_077, w_026_250, w_002_009);
  not1 I032_078(w_032_078, w_019_037);
  not1 I032_079(w_032_079, w_029_166);
  nand2 I032_081(w_032_081, w_015_034, w_017_023);
  nand2 I032_082(w_032_082, w_003_065, w_007_229);
  and2 I032_084(w_032_084, w_002_014, w_018_081);
  and2 I032_085(w_032_085, w_023_306, w_015_014);
  not1 I032_087(w_032_087, w_005_168);
  not1 I032_090(w_032_090, w_009_194);
  not1 I032_091(w_032_091, w_012_013);
  not1 I032_096(w_032_096, w_018_292);
  and2 I032_098(w_032_098, w_016_074, w_002_010);
  and2 I032_102(w_032_102, w_031_054, w_017_025);
  and2 I032_103(w_032_103, w_019_034, w_026_187);
  not1 I032_104(w_032_104, w_024_009);
  or2  I032_106(w_032_106, w_002_010, w_009_211);
  or2  I032_108(w_032_108, w_002_017, w_006_000);
  nand2 I032_110(w_032_110, w_013_106, w_022_057);
  and2 I032_114(w_032_114, w_026_386, w_029_096);
  nand2 I032_115(w_032_115, w_004_388, w_005_073);
  and2 I032_120(w_032_120, w_012_382, w_008_202);
  or2  I032_121(w_032_121, w_006_000, w_016_382);
  nand2 I032_122(w_032_122, w_021_083, w_014_065);
  and2 I032_123(w_032_123, w_009_178, w_011_106);
  and2 I032_124(w_032_124, w_016_209, w_005_172);
  or2  I032_127(w_032_127, w_022_158, w_028_395);
  and2 I032_132(w_032_132, w_029_142, w_001_004);
  nand2 I032_137(w_032_137, w_024_109, w_020_065);
  not1 I032_139(w_032_139, w_007_281);
  nand2 I032_141(w_032_141, w_010_073, w_015_134);
  not1 I032_142(w_032_142, w_020_005);
  not1 I032_143(w_032_143, w_031_014);
  and2 I032_145(w_032_145, w_027_007, w_022_132);
  not1 I032_148(w_032_148, w_005_109);
  and2 I032_153(w_032_153, w_022_099, w_029_222);
  not1 I032_154(w_032_154, w_003_006);
  or2  I032_158(w_032_158, w_015_018, w_006_000);
  not1 I032_160(w_032_160, w_007_261);
  or2  I032_165(w_032_165, w_013_039, w_025_060);
  nand2 I032_167(w_032_167, w_008_138, w_022_145);
  or2  I032_169(w_032_169, w_022_124, w_019_020);
  not1 I032_171(w_032_171, w_000_162);
  and2 I032_172(w_032_172, w_014_056, w_009_234);
  nand2 I032_176(w_032_176, w_031_050, w_018_181);
  not1 I032_177(w_032_177, w_005_216);
  and2 I032_179(w_032_179, w_002_012, w_001_001);
  or2  I032_181(w_032_181, w_005_076, w_022_088);
  and2 I032_183(w_032_183, w_024_131, w_027_027);
  or2  I032_184(w_032_184, w_015_001, w_013_123);
  nand2 I032_187(w_032_187, w_015_098, w_000_328);
  nand2 I032_188(w_032_188, w_022_105, w_030_054);
  and2 I032_190(w_032_190, w_022_158, w_029_137);
  or2  I032_195(w_032_195, w_027_035, w_013_106);
  or2  I033_000(w_033_000, w_032_049, w_000_343);
  and2 I033_001(w_033_001, w_025_104, w_005_166);
  nand2 I033_002(w_033_002, w_013_071, w_009_013);
  or2  I033_003(w_033_003, w_026_260, w_028_313);
  and2 I033_004(w_033_004, w_020_164, w_019_038);
  or2  I033_005(w_033_005, w_001_000, w_025_279);
  and2 I033_007(w_033_007, w_005_099, w_002_023);
  nand2 I033_008(w_033_008, w_016_048, w_028_011);
  or2  I033_009(w_033_009, w_020_054, w_007_060);
  not1 I033_010(w_033_010, w_006_000);
  not1 I033_011(w_033_011, w_025_105);
  and2 I033_012(w_033_012, w_024_000, w_022_049);
  or2  I033_013(w_033_013, w_002_016, w_001_004);
  and2 I033_014(w_033_014, w_007_370, w_023_325);
  or2  I033_015(w_033_015, w_006_000, w_020_154);
  not1 I033_016(w_033_016, w_008_089);
  nand2 I033_018(w_033_018, w_000_095, w_000_453);
  or2  I033_019(w_033_019, w_022_024, w_016_274);
  nand2 I033_020(w_033_020, w_017_044, w_023_058);
  not1 I033_021(w_033_021, w_011_150);
  nand2 I033_022(w_033_022, w_017_035, w_028_070);
  or2  I033_023(w_033_023, w_001_004, w_014_020);
  and2 I033_024(w_033_024, w_024_123, w_020_140);
  nand2 I033_025(w_033_025, w_018_139, w_001_006);
  not1 I033_026(w_033_026, w_017_000);
  or2  I033_027(w_033_027, w_000_428, w_028_239);
  nand2 I033_028(w_033_028, w_006_000, w_023_353);
  or2  I033_029(w_033_029, w_018_321, w_019_041);
  or2  I033_030(w_033_030, w_000_097, w_003_030);
  or2  I033_031(w_033_031, w_023_413, w_014_157);
  and2 I033_032(w_033_032, w_015_131, w_032_108);
  nand2 I033_033(w_033_033, w_006_000, w_007_231);
  or2  I033_034(w_033_034, w_023_270, w_017_033);
  nand2 I033_035(w_033_035, w_027_251, w_024_216);
  not1 I033_037(w_033_037, w_029_013);
  and2 I033_038(w_033_038, w_010_418, w_009_020);
  or2  I033_039(w_033_039, w_009_218, w_003_088);
  not1 I033_040(w_033_040, w_010_422);
  and2 I033_042(w_033_042, w_012_234, w_001_002);
  or2  I033_043(w_033_043, w_010_292, w_032_074);
  nand2 I033_044(w_033_044, w_028_335, w_021_031);
  or2  I033_045(w_033_045, w_030_027, w_029_186);
  and2 I033_046(w_033_046, w_032_181, w_026_302);
  nand2 I033_047(w_033_047, w_029_152, w_014_108);
  nand2 I033_048(w_033_048, w_024_258, w_020_180);
  not1 I033_050(w_033_050, w_027_329);
  or2  I033_051(w_033_051, w_013_091, w_020_158);
  nand2 I033_052(w_033_052, w_016_031, w_000_416);
  and2 I033_053(w_033_053, w_027_218, w_029_112);
  not1 I033_054(w_033_054, w_011_143);
  or2  I033_055(w_033_055, w_000_245, w_028_355);
  and2 I033_056(w_033_056, w_029_078, w_004_222);
  and2 I033_057(w_033_057, w_032_051, w_028_019);
  nand2 I033_058(w_033_058, w_015_092, w_010_038);
  not1 I034_003(w_034_003, w_018_001);
  or2  I034_006(w_034_006, w_005_037, w_006_000);
  or2  I034_007(w_034_007, w_016_086, w_029_014);
  nand2 I034_008(w_034_008, w_032_098, w_016_210);
  and2 I034_011(w_034_011, w_017_030, w_016_247);
  not1 I034_014(w_034_014, w_031_030);
  nand2 I034_016(w_034_016, w_021_033, w_021_005);
  or2  I034_021(w_034_021, w_021_023, w_008_300);
  and2 I034_022(w_034_022, w_006_000, w_019_030);
  and2 I034_025(w_034_025, w_028_339, w_015_095);
  or2  I034_027(w_034_027, w_014_052, w_027_018);
  not1 I034_030(w_034_030, w_014_082);
  not1 I034_031(w_034_031, w_007_167);
  and2 I034_032(w_034_032, w_003_009, w_017_023);
  nand2 I034_036(w_034_036, w_007_094, w_014_152);
  or2  I034_037(w_034_037, w_028_353, w_019_043);
  or2  I034_042(w_034_042, w_033_040, w_009_091);
  nand2 I034_043(w_034_043, w_024_093, w_024_276);
  nand2 I034_045(w_034_045, w_006_000, w_000_029);
  or2  I034_048(w_034_048, w_012_330, w_016_147);
  nand2 I034_052(w_034_052, w_026_082, w_011_039);
  and2 I034_053(w_034_053, w_032_078, w_009_147);
  and2 I034_056(w_034_056, w_019_015, w_026_022);
  not1 I034_057(w_034_057, w_030_185);
  not1 I034_058(w_034_058, w_017_191);
  and2 I034_059(w_034_059, w_012_026, w_012_094);
  and2 I034_060(w_034_060, w_033_029, w_022_121);
  nand2 I034_061(w_034_061, w_017_067, w_003_004);
  and2 I034_062(w_034_062, w_011_308, w_032_104);
  and2 I034_066(w_034_066, w_005_090, w_032_090);
  and2 I034_067(w_034_067, w_020_103, w_005_133);
  or2  I034_075(w_034_075, w_004_113, w_007_053);
  and2 I034_076(w_034_076, w_000_259, w_013_082);
  not1 I034_077(w_034_077, w_001_000);
  and2 I034_080(w_034_080, w_033_046, w_031_003);
  nand2 I034_081(w_034_081, w_010_069, w_003_054);
  not1 I034_084(w_034_084, w_029_025);
  nand2 I034_085(w_034_085, w_002_012, w_013_174);
  or2  I034_088(w_034_088, w_025_097, w_004_380);
  and2 I034_089(w_034_089, w_012_017, w_031_019);
  and2 I034_093(w_034_093, w_018_034, w_019_051);
  not1 I034_095(w_034_095, w_006_000);
  and2 I034_097(w_034_097, w_024_133, w_015_049);
  nand2 I034_098(w_034_098, w_007_176, w_029_119);
  not1 I034_100(w_034_100, w_003_019);
  or2  I034_101(w_034_101, w_030_010, w_011_292);
  nand2 I034_104(w_034_104, w_006_000, w_014_208);
  or2  I034_108(w_034_108, w_014_132, w_027_258);
  or2  I034_121(w_034_121, w_020_145, w_025_226);
  and2 I034_122(w_034_122, w_014_109, w_020_060);
  nand2 I034_124(w_034_124, w_003_044, w_013_044);
  nand2 I034_129(w_034_129, w_026_386, w_015_039);
  and2 I034_138(w_034_138, w_030_055, w_004_293);
  or2  I034_139(w_034_139, w_023_049, w_030_051);
  and2 I034_145(w_034_145, w_030_022, w_028_199);
  nand2 I034_146(w_034_146, w_025_015, w_002_009);
  not1 I034_150(w_034_150, w_019_021);
  and2 I034_152(w_034_152, w_011_339, w_004_223);
  nand2 I034_154(w_034_154, w_004_000, w_026_280);
  not1 I034_155(w_034_155, w_021_066);
  and2 I034_165(w_034_165, w_013_109, w_025_333);
  and2 I034_166(w_034_166, w_006_000, w_030_041);
  and2 I034_170(w_034_170, w_027_242, w_017_103);
  nand2 I034_172(w_034_172, w_013_062, w_023_323);
  or2  I034_177(w_034_177, w_017_181, w_015_113);
  or2  I034_179(w_034_179, w_022_101, w_024_023);
  not1 I034_182(w_034_182, w_011_296);
  and2 I034_187(w_034_187, w_029_118, w_012_345);
  and2 I034_191(w_034_191, w_003_007, w_012_366);
  not1 I034_192(w_034_192, w_028_084);
  and2 I034_193(w_034_193, w_001_001, w_014_081);
  nand2 I034_194(w_034_194, w_018_051, w_027_199);
  and2 I034_195(w_034_195, w_011_289, w_010_431);
  nand2 I034_196(w_034_196, w_031_011, w_020_033);
  or2  I034_199(w_034_199, w_024_245, w_014_165);
  nand2 I034_200(w_034_200, w_029_019, w_016_078);
  nand2 I034_202(w_034_202, w_029_067, w_014_146);
  not1 I034_203(w_034_203, w_001_006);
  and2 I034_205(w_034_205, w_012_236, w_004_016);
  or2  I034_206(w_034_206, w_003_012, w_021_038);
  and2 I034_210(w_034_210, w_025_016, w_020_043);
  or2  I034_213(w_034_213, w_000_454, w_006_000);
  and2 I034_215(w_034_215, w_009_088, w_001_004);
  and2 I034_219(w_034_219, w_024_105, w_009_000);
  not1 I034_221(w_034_221, w_001_005);
  not1 I034_222(w_034_222, w_011_188);
  nand2 I034_223(w_034_223, w_010_021, w_023_082);
  and2 I034_224(w_034_224, w_024_259, w_008_093);
  and2 I034_238(w_034_238, w_009_163, w_030_193);
  nand2 I034_240(w_034_240, w_032_071, w_026_131);
  not1 I034_247(w_034_247, w_006_000);
  not1 I034_252(w_034_252, w_032_122);
  nand2 I034_254(w_034_254, w_017_092, w_011_114);
  not1 I034_257(w_034_257, w_014_254);
  not1 I034_259(w_034_259, w_021_012);
  and2 I034_262(w_034_262, w_013_129, w_004_037);
  not1 I034_265(w_034_265, w_015_014);
  nand2 I034_267(w_034_267, w_022_069, w_024_112);
  nand2 I034_271(w_034_271, w_021_083, w_008_056);
  or2  I034_272(w_034_272, w_023_404, w_032_172);
  not1 I034_276(w_034_276, w_030_067);
  not1 I034_278(w_034_278, w_012_214);
  not1 I034_281(w_034_281, w_018_236);
  or2  I035_000(w_035_000, w_001_000, w_025_007);
  or2  I035_001(w_035_001, w_019_024, w_011_057);
  or2  I035_002(w_035_002, w_015_121, w_008_024);
  or2  I035_004(w_035_004, w_027_019, w_002_004);
  or2  I035_005(w_035_005, w_017_022, w_018_320);
  not1 I035_006(w_035_006, w_021_042);
  not1 I035_007(w_035_007, w_012_125);
  nand2 I035_008(w_035_008, w_008_027, w_013_255);
  or2  I035_009(w_035_009, w_005_228, w_007_142);
  or2  I035_010(w_035_010, w_013_109, w_020_103);
  nand2 I035_011(w_035_011, w_012_067, w_013_104);
  not1 I035_013(w_035_013, w_003_083);
  and2 I035_014(w_035_014, w_027_060, w_004_330);
  nand2 I035_015(w_035_015, w_029_189, w_001_002);
  or2  I035_016(w_035_016, w_009_213, w_002_018);
  nand2 I035_017(w_035_017, w_023_043, w_002_023);
  or2  I035_018(w_035_018, w_015_125, w_001_006);
  nand2 I035_021(w_035_021, w_013_266, w_007_072);
  or2  I035_023(w_035_023, w_024_049, w_007_173);
  not1 I035_024(w_035_024, w_022_102);
  nand2 I035_025(w_035_025, w_023_002, w_014_079);
  not1 I035_027(w_035_027, w_010_178);
  not1 I035_028(w_035_028, w_000_296);
  not1 I035_029(w_035_029, w_027_134);
  not1 I035_031(w_035_031, w_034_011);
  nand2 I035_032(w_035_032, w_034_088, w_030_160);
  nand2 I035_034(w_035_034, w_022_035, w_014_218);
  or2  I035_035(w_035_035, w_004_102, w_016_300);
  or2  I035_036(w_035_036, w_020_099, w_017_054);
  nand2 I035_037(w_035_037, w_029_217, w_027_394);
  or2  I035_038(w_035_038, w_028_005, w_011_285);
  and2 I035_039(w_035_039, w_000_312, w_012_200);
  not1 I035_040(w_035_040, w_001_005);
  not1 I035_041(w_035_041, w_027_198);
  or2  I035_045(w_035_045, w_023_016, w_032_043);
  or2  I035_046(w_035_046, w_010_159, w_020_065);
  and2 I035_047(w_035_047, w_015_078, w_015_114);
  and2 I035_048(w_035_048, w_019_002, w_029_204);
  or2  I035_049(w_035_049, w_016_122, w_024_045);
  nand2 I035_050(w_035_050, w_012_096, w_016_037);
  not1 I035_051(w_035_051, w_021_081);
  not1 I035_054(w_035_054, w_030_188);
  not1 I035_056(w_035_056, w_018_051);
  not1 I035_057(w_035_057, w_005_206);
  nand2 I035_061(w_035_061, w_021_012, w_032_115);
  nand2 I035_062(w_035_062, w_024_002, w_022_120);
  not1 I035_065(w_035_065, w_023_183);
  and2 I035_066(w_035_066, w_027_080, w_009_202);
  and2 I035_068(w_035_068, w_023_161, w_020_079);
  or2  I035_069(w_035_069, w_020_176, w_026_359);
  nand2 I035_071(w_035_071, w_003_006, w_031_034);
  nand2 I035_075(w_035_075, w_005_197, w_005_147);
  nand2 I035_077(w_035_077, w_017_007, w_003_036);
  nand2 I035_078(w_035_078, w_006_000, w_004_415);
  or2  I035_079(w_035_079, w_013_075, w_034_262);
  not1 I035_080(w_035_080, w_024_053);
  not1 I035_083(w_035_083, w_003_041);
  or2  I035_084(w_035_084, w_020_136, w_017_048);
  nand2 I035_085(w_035_085, w_000_236, w_004_278);
  not1 I035_086(w_035_086, w_029_122);
  or2  I035_088(w_035_088, w_028_008, w_008_026);
  or2  I035_089(w_035_089, w_027_088, w_013_228);
  not1 I035_090(w_035_090, w_028_325);
  nand2 I035_094(w_035_094, w_023_295, w_030_017);
  nand2 I035_096(w_035_096, w_002_003, w_031_042);
  or2  I035_097(w_035_097, w_002_007, w_005_153);
  not1 I035_100(w_035_100, w_009_133);
  or2  I035_101(w_035_101, w_017_010, w_009_067);
  nand2 I035_107(w_035_107, w_021_097, w_015_063);
  and2 I035_108(w_035_108, w_002_025, w_019_021);
  not1 I035_109(w_035_109, w_018_035);
  and2 I036_005(w_036_005, w_003_042, w_016_059);
  nand2 I036_006(w_036_006, w_022_162, w_003_001);
  nand2 I036_008(w_036_008, w_022_116, w_002_004);
  nand2 I036_016(w_036_016, w_006_000, w_004_251);
  and2 I036_017(w_036_017, w_011_112, w_001_003);
  not1 I036_025(w_036_025, w_016_328);
  nand2 I036_027(w_036_027, w_032_003, w_022_028);
  or2  I036_028(w_036_028, w_016_183, w_024_105);
  nand2 I036_030(w_036_030, w_014_007, w_007_197);
  nand2 I036_031(w_036_031, w_029_147, w_012_039);
  not1 I036_034(w_036_034, w_027_313);
  or2  I036_042(w_036_042, w_018_018, w_008_074);
  nand2 I036_043(w_036_043, w_013_180, w_027_262);
  nand2 I036_044(w_036_044, w_023_074, w_014_086);
  not1 I036_045(w_036_045, w_034_104);
  not1 I036_046(w_036_046, w_001_005);
  or2  I036_056(w_036_056, w_035_051, w_007_251);
  not1 I036_058(w_036_058, w_002_020);
  nand2 I036_060(w_036_060, w_001_005, w_020_162);
  not1 I036_061(w_036_061, w_004_216);
  nand2 I036_065(w_036_065, w_027_287, w_023_031);
  not1 I036_067(w_036_067, w_020_048);
  and2 I036_073(w_036_073, w_002_020, w_022_082);
  not1 I036_077(w_036_077, w_021_050);
  nand2 I036_078(w_036_078, w_008_020, w_032_055);
  not1 I036_079(w_036_079, w_033_003);
  not1 I036_080(w_036_080, w_035_023);
  or2  I036_081(w_036_081, w_002_018, w_032_169);
  or2  I036_084(w_036_084, w_018_083, w_021_096);
  or2  I036_087(w_036_087, w_001_003, w_018_048);
  and2 I036_093(w_036_093, w_023_374, w_025_261);
  or2  I036_094(w_036_094, w_020_096, w_005_101);
  and2 I036_095(w_036_095, w_023_068, w_014_091);
  nand2 I036_098(w_036_098, w_034_221, w_029_176);
  not1 I036_099(w_036_099, w_017_115);
  nand2 I036_101(w_036_101, w_031_024, w_007_029);
  or2  I036_105(w_036_105, w_023_061, w_019_032);
  not1 I036_108(w_036_108, w_000_036);
  or2  I036_113(w_036_113, w_021_026, w_001_001);
  and2 I036_118(w_036_118, w_017_104, w_001_001);
  or2  I036_120(w_036_120, w_029_124, w_008_140);
  not1 I036_127(w_036_127, w_015_059);
  not1 I036_128(w_036_128, w_001_001);
  or2  I036_129(w_036_129, w_004_010, w_029_141);
  or2  I036_131(w_036_131, w_027_031, w_020_071);
  and2 I036_141(w_036_141, w_008_070, w_035_025);
  nand2 I036_143(w_036_143, w_018_249, w_031_020);
  or2  I036_147(w_036_147, w_032_184, w_005_143);
  not1 I036_152(w_036_152, w_015_121);
  not1 I036_155(w_036_155, w_013_255);
  not1 I036_157(w_036_157, w_005_022);
  nand2 I036_163(w_036_163, w_030_113, w_022_116);
  not1 I036_165(w_036_165, w_024_211);
  and2 I036_166(w_036_166, w_002_024, w_025_413);
  nand2 I036_168(w_036_168, w_028_035, w_000_075);
  not1 I036_169(w_036_169, w_027_268);
  not1 I036_171(w_036_171, w_030_078);
  and2 I036_175(w_036_175, w_022_009, w_016_099);
  and2 I036_179(w_036_179, w_008_242, w_006_000);
  and2 I036_181(w_036_181, w_021_059, w_006_000);
  or2  I036_184(w_036_184, w_018_000, w_011_153);
  or2  I036_188(w_036_188, w_023_271, w_020_159);
  not1 I036_190(w_036_190, w_030_090);
  and2 I036_195(w_036_195, w_012_061, w_000_236);
  and2 I036_196(w_036_196, w_009_175, w_029_121);
  not1 I036_200(w_036_200, w_028_087);
  or2  I036_201(w_036_201, w_025_450, w_025_420);
  nand2 I036_202(w_036_202, w_012_348, w_008_177);
  nand2 I036_204(w_036_204, w_022_118, w_027_153);
  and2 I036_205(w_036_205, w_011_061, w_031_004);
  not1 I036_209(w_036_209, w_005_113);
  and2 I036_216(w_036_216, w_035_049, w_033_033);
  nand2 I036_219(w_036_219, w_024_070, w_006_000);
  and2 I036_227(w_036_227, w_035_062, w_017_033);
  nand2 I036_229(w_036_229, w_016_022, w_027_011);
  or2  I036_234(w_036_234, w_019_006, w_016_347);
  nand2 I036_260(w_036_260, w_003_096, w_033_042);
  and2 I036_261(w_036_261, w_016_077, w_004_065);
  and2 I036_272(w_036_272, w_009_197, w_012_174);
  and2 I036_278(w_036_278, w_017_081, w_019_040);
  nand2 I037_001(w_037_001, w_009_213, w_009_223);
  nand2 I037_002(w_037_002, w_024_087, w_029_231);
  not1 I037_004(w_037_004, w_002_013);
  not1 I037_010(w_037_010, w_020_048);
  and2 I037_011(w_037_011, w_015_106, w_036_017);
  and2 I037_013(w_037_013, w_020_186, w_008_186);
  nand2 I037_014(w_037_014, w_029_192, w_022_002);
  not1 I037_015(w_037_015, w_027_022);
  not1 I037_018(w_037_018, w_019_015);
  not1 I037_020(w_037_020, w_023_311);
  not1 I037_021(w_037_021, w_021_042);
  nand2 I037_022(w_037_022, w_006_000, w_020_183);
  not1 I037_023(w_037_023, w_025_477);
  nand2 I037_024(w_037_024, w_034_006, w_007_239);
  not1 I037_029(w_037_029, w_034_215);
  not1 I037_030(w_037_030, w_000_455);
  nand2 I037_031(w_037_031, w_026_342, w_021_000);
  not1 I037_032(w_037_032, w_003_084);
  or2  I037_035(w_037_035, w_028_009, w_023_191);
  or2  I037_036(w_037_036, w_009_130, w_013_005);
  not1 I037_037(w_037_037, w_032_084);
  and2 I037_038(w_037_038, w_024_143, w_035_025);
  and2 I037_041(w_037_041, w_021_060, w_018_229);
  nand2 I037_042(w_037_042, w_004_272, w_023_145);
  nand2 I037_043(w_037_043, w_014_151, w_032_120);
  nand2 I037_047(w_037_047, w_032_053, w_019_024);
  or2  I037_048(w_037_048, w_000_375, w_013_113);
  nand2 I037_049(w_037_049, w_014_027, w_020_011);
  not1 I037_050(w_037_050, w_030_118);
  or2  I037_052(w_037_052, w_015_001, w_025_428);
  nand2 I037_053(w_037_053, w_022_140, w_014_114);
  or2  I037_057(w_037_057, w_003_086, w_028_241);
  and2 I037_058(w_037_058, w_009_212, w_007_087);
  nand2 I037_059(w_037_059, w_011_272, w_020_186);
  not1 I037_060(w_037_060, w_012_300);
  nand2 I037_064(w_037_064, w_018_084, w_008_237);
  nand2 I037_065(w_037_065, w_002_009, w_024_133);
  not1 I037_066(w_037_066, w_026_021);
  and2 I037_067(w_037_067, w_003_045, w_015_116);
  nand2 I037_068(w_037_068, w_022_051, w_006_000);
  or2  I037_069(w_037_069, w_018_131, w_020_019);
  or2  I037_072(w_037_072, w_020_083, w_025_233);
  not1 I037_075(w_037_075, w_031_066);
  not1 I037_076(w_037_076, w_029_006);
  and2 I037_078(w_037_078, w_033_057, w_014_080);
  and2 I037_081(w_037_081, w_022_154, w_004_431);
  or2  I037_084(w_037_084, w_018_248, w_027_063);
  or2  I037_085(w_037_085, w_019_035, w_017_071);
  nand2 I037_086(w_037_086, w_010_170, w_030_006);
  or2  I037_087(w_037_087, w_005_217, w_012_294);
  and2 I037_089(w_037_089, w_029_163, w_031_021);
  not1 I037_090(w_037_090, w_019_004);
  not1 I037_091(w_037_091, w_009_181);
  not1 I037_093(w_037_093, w_015_024);
  and2 I037_097(w_037_097, w_023_196, w_004_144);
  and2 I037_100(w_037_100, w_001_005, w_032_121);
  not1 I037_101(w_037_101, w_014_231);
  and2 I037_114(w_037_114, w_034_199, w_027_039);
  or2  I037_115(w_037_115, w_034_259, w_009_186);
  not1 I037_116(w_037_116, w_009_206);
  or2  I037_117(w_037_117, w_021_024, w_003_036);
  or2  I037_118(w_037_118, w_035_077, w_009_083);
  and2 I037_119(w_037_119, w_015_000, w_012_071);
  or2  I037_120(w_037_120, w_007_262, w_004_260);
  or2  I037_121(w_037_121, w_031_027, w_024_037);
  not1 I037_122(w_037_122, w_011_033);
  nand2 I037_124(w_037_124, w_027_412, w_006_000);
  and2 I037_125(w_037_125, w_030_124, w_032_143);
  and2 I037_126(w_037_126, w_007_045, w_025_094);
  and2 I037_127(w_037_127, w_029_107, w_012_122);
  not1 I037_128(w_037_128, w_014_047);
  and2 I037_130(w_037_130, w_036_093, w_009_232);
  not1 I037_132(w_037_132, w_024_186);
  or2  I037_138(w_037_138, w_008_091, w_000_065);
  or2  I037_140(w_037_140, w_005_103, w_002_014);
  nand2 I037_142(w_037_142, w_034_098, w_007_403);
  not1 I037_143(w_037_143, w_036_079);
  not1 I037_144(w_037_144, w_019_033);
  or2  I037_149(w_037_149, w_021_041, w_000_457);
  and2 I038_000(w_038_000, w_031_033, w_004_228);
  and2 I038_001(w_038_001, w_008_102, w_011_242);
  nand2 I038_002(w_038_002, w_032_123, w_008_064);
  nand2 I038_005(w_038_005, w_012_028, w_003_068);
  and2 I038_007(w_038_007, w_020_053, w_031_019);
  not1 I038_008(w_038_008, w_014_039);
  or2  I038_009(w_038_009, w_000_222, w_004_085);
  not1 I038_010(w_038_010, w_000_401);
  nand2 I038_011(w_038_011, w_012_080, w_003_094);
  not1 I038_012(w_038_012, w_015_088);
  not1 I038_013(w_038_013, w_014_044);
  not1 I038_014(w_038_014, w_022_090);
  not1 I038_016(w_038_016, w_015_063);
  and2 I038_019(w_038_019, w_037_058, w_014_183);
  or2  I038_020(w_038_020, w_033_025, w_023_006);
  not1 I038_021(w_038_021, w_025_130);
  not1 I038_022(w_038_022, w_037_142);
  and2 I038_023(w_038_023, w_035_077, w_034_108);
  not1 I038_024(w_038_024, w_033_047);
  not1 I038_026(w_038_026, w_006_000);
  not1 I038_028(w_038_028, w_030_047);
  and2 I038_030(w_038_030, w_029_231, w_005_176);
  and2 I038_031(w_038_031, w_001_002, w_011_115);
  nand2 I038_032(w_038_032, w_025_012, w_008_124);
  and2 I038_035(w_038_035, w_000_452, w_016_189);
  nand2 I038_037(w_038_037, w_020_131, w_016_022);
  and2 I038_040(w_038_040, w_002_020, w_026_341);
  or2  I038_041(w_038_041, w_024_044, w_023_165);
  and2 I038_044(w_038_044, w_007_359, w_020_107);
  and2 I038_046(w_038_046, w_026_014, w_008_035);
  and2 I038_047(w_038_047, w_008_125, w_021_035);
  and2 I038_049(w_038_049, w_006_000, w_010_181);
  or2  I038_051(w_038_051, w_018_091, w_013_068);
  not1 I038_054(w_038_054, w_023_210);
  and2 I038_055(w_038_055, w_033_022, w_032_190);
  not1 I038_056(w_038_056, w_021_086);
  and2 I038_058(w_038_058, w_026_367, w_005_108);
  or2  I038_062(w_038_062, w_012_006, w_017_018);
  or2  I038_064(w_038_064, w_022_121, w_025_095);
  and2 I038_066(w_038_066, w_035_001, w_025_349);
  nand2 I038_067(w_038_067, w_032_026, w_015_068);
  not1 I038_068(w_038_068, w_020_091);
  and2 I038_069(w_038_069, w_037_038, w_035_032);
  and2 I038_070(w_038_070, w_037_084, w_010_197);
  nand2 I038_073(w_038_073, w_011_220, w_032_054);
  nand2 I038_074(w_038_074, w_004_472, w_016_330);
  nand2 I038_075(w_038_075, w_014_108, w_009_200);
  and2 I038_077(w_038_077, w_033_038, w_006_000);
  nand2 I038_079(w_038_079, w_022_127, w_029_172);
  or2  I038_080(w_038_080, w_009_163, w_001_005);
  or2  I038_081(w_038_081, w_036_042, w_036_128);
  not1 I038_082(w_038_082, w_000_458);
  or2  I038_086(w_038_086, w_012_356, w_028_049);
  nand2 I038_087(w_038_087, w_036_171, w_003_005);
  not1 I038_088(w_038_088, w_018_123);
  or2  I038_089(w_038_089, w_000_263, w_007_106);
  nand2 I038_093(w_038_093, w_021_093, w_036_108);
  and2 I038_094(w_038_094, w_017_065, w_016_268);
  not1 I038_096(w_038_096, w_029_213);
  or2  I038_099(w_038_099, w_005_179, w_000_411);
  nand2 I039_001(w_039_001, w_000_433, w_022_046);
  not1 I039_002(w_039_002, w_012_020);
  nand2 I039_014(w_039_014, w_006_000, w_035_002);
  or2  I039_024(w_039_024, w_001_006, w_029_136);
  or2  I039_040(w_039_040, w_036_278, w_010_115);
  or2  I039_046(w_039_046, w_034_030, w_029_045);
  nand2 I039_048(w_039_048, w_030_090, w_002_024);
  not1 I039_056(w_039_056, w_024_122);
  or2  I039_057(w_039_057, w_025_113, w_021_073);
  not1 I039_060(w_039_060, w_014_225);
  or2  I039_063(w_039_063, w_008_078, w_006_000);
  not1 I039_067(w_039_067, w_024_185);
  not1 I039_077(w_039_077, w_005_037);
  not1 I039_080(w_039_080, w_005_104);
  not1 I039_083(w_039_083, w_032_148);
  and2 I039_085(w_039_085, w_032_015, w_008_198);
  or2  I039_089(w_039_089, w_030_097, w_020_023);
  or2  I039_093(w_039_093, w_008_060, w_031_010);
  and2 I039_100(w_039_100, w_015_121, w_001_004);
  nand2 I039_103(w_039_103, w_014_065, w_013_011);
  and2 I039_104(w_039_104, w_028_039, w_026_341);
  not1 I039_107(w_039_107, w_027_240);
  and2 I039_108(w_039_108, w_013_044, w_031_045);
  not1 I039_109(w_039_109, w_022_038);
  not1 I039_111(w_039_111, w_025_143);
  and2 I039_113(w_039_113, w_001_004, w_010_361);
  not1 I039_117(w_039_117, w_003_042);
  not1 I039_130(w_039_130, w_016_399);
  or2  I039_136(w_039_136, w_009_032, w_032_181);
  nand2 I039_145(w_039_145, w_017_173, w_006_000);
  and2 I039_146(w_039_146, w_005_078, w_015_005);
  nand2 I039_151(w_039_151, w_003_041, w_002_013);
  or2  I039_153(w_039_153, w_003_007, w_029_178);
  and2 I039_158(w_039_158, w_004_385, w_023_318);
  nand2 I039_160(w_039_160, w_007_349, w_019_028);
  not1 I039_176(w_039_176, w_000_064);
  not1 I039_177(w_039_177, w_023_058);
  and2 I039_182(w_039_182, w_014_249, w_000_141);
  and2 I039_191(w_039_191, w_029_151, w_008_064);
  not1 I039_198(w_039_198, w_013_118);
  and2 I039_204(w_039_204, w_038_000, w_027_112);
  or2  I039_212(w_039_212, w_012_101, w_034_265);
  not1 I039_215(w_039_215, w_006_000);
  or2  I039_216(w_039_216, w_026_148, w_000_380);
  not1 I039_220(w_039_220, w_012_258);
  nand2 I039_221(w_039_221, w_025_429, w_016_301);
  and2 I039_223(w_039_223, w_020_003, w_026_375);
  nand2 I039_224(w_039_224, w_033_048, w_006_000);
  nand2 I039_225(w_039_225, w_005_179, w_026_012);
  not1 I039_237(w_039_237, w_004_010);
  not1 I039_240(w_039_240, w_011_099);
  not1 I039_241(w_039_241, w_019_037);
  and2 I039_250(w_039_250, w_000_014, w_034_104);
  and2 I039_254(w_039_254, w_034_007, w_031_000);
  not1 I039_268(w_039_268, w_007_302);
  not1 I039_270(w_039_270, w_033_022);
  or2  I039_272(w_039_272, w_036_084, w_007_006);
  and2 I039_274(w_039_274, w_017_086, w_027_141);
  and2 I039_278(w_039_278, w_002_027, w_034_095);
  not1 I039_292(w_039_292, w_014_040);
  and2 I039_295(w_039_295, w_009_104, w_033_007);
  not1 I039_306(w_039_306, w_038_082);
  not1 I039_309(w_039_309, w_009_109);
  or2  I039_331(w_039_331, w_017_000, w_013_218);
  not1 I039_334(w_039_334, w_015_071);
  nand2 I039_337(w_039_337, w_030_081, w_036_195);
  not1 I039_338(w_039_338, w_003_007);
  or2  I039_343(w_039_343, w_005_239, w_024_191);
  not1 I039_344(w_039_344, w_004_125);
  nand2 I039_346(w_039_346, w_028_014, w_009_222);
  and2 I039_348(w_039_348, w_006_000, w_036_165);
  or2  I039_354(w_039_354, w_013_155, w_003_033);
  or2  I039_356(w_039_356, w_023_038, w_011_099);
  not1 I039_357(w_039_357, w_031_029);
  not1 I039_364(w_039_364, w_028_035);
  nand2 I039_366(w_039_366, w_001_000, w_030_119);
  and2 I039_367(w_039_367, w_014_195, w_017_019);
  nand2 I039_370(w_039_370, w_008_193, w_027_366);
  or2  I039_374(w_039_374, w_018_146, w_005_053);
  not1 I039_376(w_039_376, w_001_003);
  nand2 I039_381(w_039_381, w_030_119, w_006_000);
  and2 I039_394(w_039_394, w_007_284, w_009_206);
  and2 I039_395(w_039_395, w_022_101, w_012_026);
  or2  I039_396(w_039_396, w_023_010, w_002_020);
  not1 I039_397(w_039_397, w_002_015);
  nand2 I039_400(w_039_400, w_017_141, w_014_247);
  and2 I039_402(w_039_402, w_005_181, w_009_223);
  nand2 I039_404(w_039_404, w_033_051, w_022_122);
  and2 I039_421(w_039_421, w_034_016, w_033_026);
  or2  I039_435(w_039_435, w_026_316, w_032_013);
  nand2 I039_441(w_039_441, w_009_127, w_038_046);
  not1 I039_448(w_039_448, w_001_003);
  and2 I039_451(w_039_451, w_033_027, w_006_000);
  not1 I039_454(w_039_454, w_024_096);
  not1 I039_463(w_039_463, w_015_115);
  and2 I039_475(w_039_475, w_027_169, w_000_455);
  or2  I039_483(w_039_483, w_019_012, w_011_340);
  not1 I039_494(w_039_494, w_038_049);
  not1 I039_496(w_039_496, w_008_105);
  or2  I039_498(w_039_500, w_039_499, w_039_522);
  and2 I039_499(w_039_501, w_039_500, w_035_031);
  nand2 I039_500(w_039_502, w_039_501, w_007_281);
  and2 I039_501(w_039_503, w_013_022, w_039_502);
  or2  I039_502(w_039_504, w_034_138, w_039_503);
  not1 I039_503(w_039_505, w_039_504);
  or2  I039_504(w_039_506, w_039_505, w_019_017);
  nand2 I039_505(w_039_507, w_027_217, w_039_506);
  not1 I039_506(w_039_508, w_039_507);
  not1 I039_507(w_039_509, w_039_508);
  nand2 I039_508(w_039_499, w_003_015, w_039_509);
  not1 I039_509(w_039_514, w_039_513);
  or2  I039_510(w_039_515, w_034_022, w_039_514);
  not1 I039_511(w_039_516, w_039_515);
  or2  I039_512(w_039_517, w_039_516, w_033_018);
  nand2 I039_513(w_039_518, w_039_517, w_035_035);
  and2 I039_514(w_039_519, w_003_078, w_039_518);
  not1 I039_515(w_039_520, w_039_519);
  not1 I039_516(w_039_513, w_039_500);
  and2 I039_517(w_039_522, w_037_035, w_039_520);
  and2 I040_000(w_040_000, w_031_011, w_024_046);
  nand2 I040_001(w_040_001, w_021_076, w_008_065);
  not1 I040_002(w_040_002, w_020_089);
  and2 I040_003(w_040_003, w_034_276, w_016_003);
  or2  I040_004(w_040_004, w_015_014, w_018_030);
  not1 I040_005(w_040_005, w_029_149);
  and2 I040_006(w_040_006, w_016_391, w_014_024);
  or2  I041_000(w_041_000, w_029_059, w_039_158);
  and2 I041_003(w_041_003, w_007_259, w_030_157);
  not1 I041_004(w_041_004, w_004_255);
  or2  I041_006(w_041_006, w_040_000, w_000_448);
  nand2 I041_007(w_041_007, w_031_008, w_034_222);
  nand2 I041_011(w_041_011, w_008_016, w_019_040);
  or2  I041_013(w_041_013, w_036_025, w_034_152);
  nand2 I041_022(w_041_022, w_000_275, w_038_067);
  or2  I041_024(w_041_024, w_036_204, w_025_396);
  or2  I041_025(w_041_025, w_010_338, w_039_103);
  nand2 I041_031(w_041_031, w_022_106, w_021_001);
  and2 I041_033(w_041_033, w_013_175, w_004_152);
  not1 I041_036(w_041_036, w_006_000);
  not1 I041_037(w_041_037, w_016_244);
  not1 I041_038(w_041_038, w_012_091);
  nand2 I041_039(w_041_039, w_019_007, w_033_056);
  nand2 I041_040(w_041_040, w_003_060, w_035_032);
  nand2 I041_048(w_041_048, w_012_043, w_026_060);
  or2  I041_052(w_041_052, w_010_322, w_036_101);
  and2 I041_056(w_041_056, w_038_007, w_003_035);
  not1 I041_058(w_041_058, w_007_215);
  nand2 I041_059(w_041_059, w_020_016, w_031_004);
  nand2 I041_064(w_041_064, w_035_021, w_020_155);
  nand2 I041_065(w_041_065, w_028_058, w_025_137);
  and2 I041_071(w_041_071, w_028_151, w_003_039);
  or2  I041_072(w_041_072, w_030_180, w_022_157);
  or2  I041_073(w_041_073, w_008_033, w_007_080);
  not1 I041_075(w_041_075, w_007_227);
  not1 I041_077(w_041_077, w_028_060);
  or2  I041_081(w_041_081, w_029_121, w_021_072);
  not1 I041_087(w_041_087, w_006_000);
  nand2 I041_088(w_041_088, w_035_054, w_004_340);
  nand2 I041_091(w_041_091, w_002_027, w_006_000);
  and2 I041_096(w_041_096, w_001_005, w_017_155);
  or2  I041_098(w_041_098, w_037_024, w_006_000);
  not1 I041_099(w_041_099, w_022_123);
  and2 I041_101(w_041_101, w_031_040, w_037_100);
  nand2 I041_109(w_041_109, w_025_404, w_014_153);
  and2 I041_113(w_041_113, w_000_323, w_033_012);
  nand2 I041_114(w_041_114, w_022_115, w_019_015);
  and2 I041_122(w_041_122, w_011_327, w_008_258);
  nand2 I041_125(w_041_125, w_034_045, w_036_065);
  not1 I041_128(w_041_128, w_019_000);
  nand2 I041_129(w_041_129, w_005_245, w_007_354);
  or2  I041_130(w_041_130, w_000_163, w_001_005);
  and2 I041_132(w_041_132, w_002_017, w_031_067);
  not1 I041_135(w_041_135, w_020_059);
  or2  I041_136(w_041_136, w_025_030, w_024_061);
  and2 I041_138(w_041_138, w_023_395, w_021_066);
  nand2 I041_139(w_041_139, w_026_087, w_034_165);
  or2  I041_140(w_041_140, w_024_109, w_002_006);
  or2  I041_141(w_041_141, w_001_002, w_016_255);
  nand2 I041_142(w_041_142, w_033_050, w_015_045);
  and2 I041_147(w_041_147, w_026_201, w_022_141);
  and2 I041_150(w_041_150, w_033_008, w_025_422);
  or2  I041_151(w_041_151, w_040_002, w_010_326);
  not1 I041_154(w_041_154, w_001_001);
  not1 I041_155(w_041_155, w_031_051);
  not1 I041_160(w_041_160, w_040_001);
  and2 I041_164(w_041_164, w_038_028, w_009_101);
  nand2 I041_167(w_041_167, w_019_053, w_023_270);
  not1 I041_168(w_041_168, w_007_088);
  not1 I041_169(w_041_169, w_037_101);
  not1 I041_173(w_041_173, w_008_280);
  and2 I041_175(w_041_175, w_022_146, w_008_086);
  not1 I041_182(w_041_182, w_031_056);
  not1 I041_185(w_041_185, w_038_069);
  nand2 I041_186(w_041_186, w_031_046, w_035_010);
  not1 I041_195(w_041_195, w_037_090);
  not1 I041_207(w_041_207, w_020_124);
  and2 I041_208(w_041_208, w_035_050, w_014_048);
  or2  I041_211(w_041_211, w_020_020, w_007_170);
  and2 I041_214(w_041_214, w_005_156, w_002_010);
  and2 I041_217(w_041_217, w_038_094, w_037_035);
  not1 I041_222(w_041_222, w_024_036);
  or2  I041_223(w_041_223, w_039_366, w_005_085);
  and2 I041_228(w_041_228, w_023_348, w_000_352);
  nand2 I041_235(w_041_235, w_008_324, w_007_159);
  nand2 I041_241(w_041_241, w_032_002, w_015_029);
  nand2 I041_255(w_041_255, w_026_014, w_000_091);
  and2 I041_260(w_041_260, w_005_031, w_005_246);
  not1 I041_271(w_041_271, w_026_011);
  and2 I041_288(w_041_288, w_013_001, w_007_356);
  nand2 I041_291(w_041_291, w_003_044, w_040_003);
  nand2 I041_295(w_041_295, w_002_012, w_020_101);
  not1 I041_298(w_041_298, w_007_075);
  not1 I041_300(w_041_300, w_028_085);
  nand2 I042_001(w_042_001, w_004_449, w_023_218);
  nand2 I042_002(w_042_002, w_012_050, w_004_154);
  nand2 I042_005(w_042_005, w_030_035, w_028_324);
  and2 I042_013(w_042_013, w_028_305, w_018_250);
  not1 I042_016(w_042_016, w_013_268);
  nand2 I042_033(w_042_033, w_030_019, w_010_254);
  nand2 I042_040(w_042_040, w_010_443, w_030_186);
  or2  I042_044(w_042_044, w_000_462, w_038_010);
  not1 I042_047(w_042_047, w_012_197);
  or2  I042_051(w_042_051, w_012_184, w_034_121);
  nand2 I042_054(w_042_054, w_014_155, w_032_084);
  and2 I042_055(w_042_055, w_041_136, w_010_180);
  or2  I042_058(w_042_058, w_001_000, w_036_163);
  nand2 I042_065(w_042_065, w_002_004, w_033_046);
  nand2 I042_067(w_042_067, w_035_075, w_025_470);
  or2  I042_072(w_042_072, w_034_060, w_001_006);
  nand2 I042_073(w_042_073, w_038_035, w_016_017);
  and2 I042_075(w_042_075, w_029_061, w_013_201);
  not1 I042_077(w_042_077, w_023_325);
  not1 I042_078(w_042_078, w_008_087);
  nand2 I042_082(w_042_082, w_036_196, w_008_161);
  or2  I042_084(w_042_084, w_024_163, w_000_213);
  nand2 I042_088(w_042_088, w_017_028, w_019_000);
  or2  I042_092(w_042_092, w_033_046, w_026_142);
  and2 I042_094(w_042_094, w_010_406, w_030_022);
  and2 I042_096(w_042_096, w_022_133, w_009_196);
  nand2 I042_099(w_042_099, w_023_401, w_020_046);
  or2  I042_101(w_042_101, w_002_007, w_029_017);
  or2  I042_102(w_042_102, w_003_027, w_035_028);
  and2 I042_106(w_042_106, w_032_167, w_008_212);
  or2  I042_108(w_042_108, w_000_198, w_005_038);
  and2 I042_110(w_042_110, w_025_009, w_030_172);
  not1 I042_111(w_042_111, w_026_133);
  and2 I042_113(w_042_113, w_009_132, w_000_339);
  or2  I042_120(w_042_120, w_005_232, w_010_268);
  or2  I042_121(w_042_121, w_000_104, w_025_463);
  not1 I042_126(w_042_126, w_005_126);
  or2  I042_131(w_042_131, w_038_064, w_014_035);
  nand2 I042_133(w_042_133, w_035_035, w_014_227);
  not1 I042_134(w_042_134, w_024_100);
  and2 I042_138(w_042_138, w_028_335, w_036_073);
  and2 I042_142(w_042_142, w_041_072, w_024_052);
  or2  I042_145(w_042_145, w_027_263, w_008_047);
  and2 I042_152(w_042_152, w_027_403, w_006_000);
  not1 I042_154(w_042_154, w_034_213);
  nand2 I042_158(w_042_158, w_041_122, w_018_118);
  and2 I042_160(w_042_160, w_026_387, w_014_122);
  nand2 I042_163(w_042_163, w_027_452, w_008_287);
  or2  I042_166(w_042_166, w_020_145, w_039_496);
  nand2 I042_169(w_042_169, w_037_021, w_023_251);
  and2 I042_170(w_042_170, w_022_131, w_029_221);
  nand2 I042_177(w_042_177, w_039_292, w_013_189);
  nand2 I042_178(w_042_178, w_030_043, w_032_078);
  and2 I042_183(w_042_183, w_020_186, w_013_160);
  nand2 I042_187(w_042_187, w_030_031, w_021_032);
  not1 I042_188(w_042_188, w_010_038);
  or2  I042_189(w_042_189, w_038_088, w_026_180);
  and2 I042_193(w_042_193, w_000_463, w_005_141);
  and2 I042_196(w_042_196, w_008_076, w_022_036);
  not1 I042_199(w_042_199, w_018_199);
  not1 I042_200(w_042_200, w_019_049);
  or2  I042_202(w_042_202, w_022_098, w_019_013);
  and2 I042_206(w_042_206, w_008_218, w_036_201);
  or2  I042_212(w_042_212, w_041_128, w_006_000);
  and2 I042_217(w_042_217, w_034_052, w_012_187);
  nand2 I042_221(w_042_221, w_015_080, w_032_053);
  nand2 I042_223(w_042_223, w_019_030, w_041_298);
  not1 I042_232(w_042_232, w_024_049);
  or2  I042_234(w_042_234, w_006_000, w_018_032);
  nand2 I042_250(w_042_250, w_040_000, w_013_020);
  and2 I042_255(w_042_255, w_010_121, w_021_088);
  or2  I042_265(w_042_265, w_021_091, w_008_216);
  and2 I042_270(w_042_270, w_024_179, w_040_006);
  or2  I042_275(w_042_275, w_028_381, w_003_069);
  nand2 I043_000(w_043_000, w_019_025, w_028_042);
  nand2 I043_006(w_043_006, w_026_342, w_028_208);
  and2 I043_007(w_043_007, w_019_008, w_024_009);
  or2  I043_011(w_043_011, w_035_001, w_026_332);
  not1 I043_014(w_043_014, w_016_182);
  and2 I043_016(w_043_016, w_007_125, w_029_157);
  and2 I043_019(w_043_019, w_022_003, w_029_099);
  or2  I043_022(w_043_022, w_002_011, w_008_070);
  or2  I043_026(w_043_026, w_013_117, w_020_167);
  and2 I043_029(w_043_029, w_026_377, w_033_010);
  nand2 I043_032(w_043_032, w_009_083, w_010_377);
  or2  I043_035(w_043_035, w_007_329, w_027_178);
  not1 I043_037(w_043_037, w_034_025);
  not1 I043_043(w_043_043, w_011_051);
  nand2 I043_052(w_043_052, w_032_096, w_000_276);
  and2 I043_056(w_043_056, w_009_228, w_017_081);
  and2 I043_059(w_043_059, w_022_161, w_009_038);
  or2  I043_060(w_043_060, w_010_053, w_011_018);
  and2 I043_063(w_043_063, w_037_118, w_028_236);
  not1 I043_064(w_043_064, w_015_038);
  or2  I043_065(w_043_065, w_040_001, w_020_138);
  or2  I043_069(w_043_069, w_011_136, w_027_328);
  and2 I043_071(w_043_071, w_020_039, w_037_138);
  or2  I043_077(w_043_077, w_027_166, w_018_040);
  nand2 I043_080(w_043_080, w_006_000, w_013_250);
  or2  I043_082(w_043_082, w_038_066, w_027_367);
  nand2 I043_089(w_043_089, w_030_160, w_013_144);
  nand2 I043_092(w_043_092, w_008_054, w_034_206);
  or2  I043_093(w_043_093, w_000_284, w_008_038);
  nand2 I043_094(w_043_094, w_031_013, w_027_150);
  or2  I043_099(w_043_099, w_025_014, w_041_182);
  not1 I043_101(w_043_101, w_026_150);
  and2 I043_103(w_043_103, w_036_216, w_006_000);
  or2  I043_111(w_043_111, w_027_032, w_032_114);
  not1 I043_113(w_043_113, w_011_077);
  not1 I043_119(w_043_119, w_013_035);
  nand2 I043_121(w_043_121, w_021_090, w_002_004);
  not1 I043_129(w_043_129, w_033_042);
  not1 I043_139(w_043_139, w_023_231);
  not1 I043_141(w_043_141, w_001_004);
  nand2 I043_143(w_043_143, w_017_109, w_022_035);
  nand2 I043_156(w_043_156, w_027_067, w_033_009);
  and2 I043_161(w_043_161, w_030_035, w_019_021);
  not1 I043_171(w_043_171, w_036_129);
  nand2 I043_174(w_043_174, w_028_335, w_017_043);
  not1 I043_179(w_043_179, w_005_050);
  or2  I043_183(w_043_183, w_040_005, w_020_139);
  nand2 I043_190(w_043_190, w_003_086, w_021_020);
  and2 I043_192(w_043_192, w_018_211, w_031_012);
  nand2 I043_198(w_043_198, w_018_151, w_014_152);
  nand2 I043_202(w_043_202, w_002_016, w_028_108);
  not1 I043_206(w_043_206, w_028_296);
  or2  I043_211(w_043_211, w_032_079, w_022_000);
  not1 I043_212(w_043_212, w_035_036);
  or2  I043_215(w_043_215, w_016_152, w_011_187);
  nand2 I043_217(w_043_217, w_034_053, w_007_362);
  nand2 I043_218(w_043_218, w_039_441, w_015_012);
  or2  I043_222(w_043_222, w_040_004, w_016_234);
  and2 I043_225(w_043_225, w_014_159, w_040_004);
  nand2 I043_226(w_043_226, w_005_025, w_013_204);
  not1 I043_227(w_043_227, w_028_016);
  not1 I043_230(w_043_230, w_029_080);
  and2 I043_233(w_043_233, w_031_031, w_008_011);
  nand2 I043_237(w_043_237, w_006_000, w_011_296);
  nand2 I043_238(w_043_238, w_019_044, w_021_099);
  or2  I043_241(w_043_241, w_034_056, w_006_000);
  and2 I043_242(w_043_242, w_016_187, w_014_265);
  and2 I044_001(w_044_001, w_040_006, w_043_035);
  or2  I044_007(w_044_007, w_001_003, w_040_004);
  nand2 I044_008(w_044_008, w_013_149, w_006_000);
  or2  I044_013(w_044_013, w_030_040, w_039_191);
  nand2 I044_014(w_044_014, w_011_334, w_014_102);
  or2  I044_018(w_044_018, w_032_035, w_012_364);
  and2 I044_021(w_044_021, w_033_005, w_036_202);
  or2  I044_023(w_044_023, w_041_040, w_043_111);
  and2 I044_025(w_044_025, w_003_053, w_028_341);
  and2 I044_028(w_044_028, w_031_010, w_042_082);
  nand2 I044_032(w_044_032, w_005_041, w_033_045);
  and2 I044_034(w_044_034, w_032_165, w_040_003);
  or2  I044_036(w_044_036, w_010_322, w_016_125);
  and2 I044_037(w_044_037, w_012_116, w_041_073);
  or2  I044_038(w_044_038, w_037_048, w_040_004);
  nand2 I044_048(w_044_048, w_011_018, w_011_027);
  not1 I044_049(w_044_049, w_000_055);
  not1 I044_050(w_044_050, w_006_000);
  or2  I044_053(w_044_053, w_035_089, w_014_027);
  or2  I044_055(w_044_055, w_025_260, w_040_002);
  or2  I044_059(w_044_059, w_001_001, w_006_000);
  nand2 I044_062(w_044_062, w_012_314, w_018_119);
  not1 I044_070(w_044_070, w_029_029);
  or2  I044_073(w_044_073, w_022_074, w_003_024);
  not1 I044_074(w_044_074, w_005_058);
  nand2 I044_075(w_044_075, w_016_355, w_015_005);
  and2 I044_087(w_044_087, w_030_006, w_028_309);
  not1 I044_091(w_044_091, w_035_045);
  and2 I044_094(w_044_094, w_021_094, w_030_056);
  or2  I044_101(w_044_101, w_039_117, w_040_005);
  and2 I044_108(w_044_108, w_025_127, w_003_047);
  not1 I044_109(w_044_109, w_027_370);
  nand2 I044_110(w_044_110, w_024_250, w_039_089);
  nand2 I044_112(w_044_112, w_010_398, w_000_125);
  nand2 I044_119(w_044_119, w_039_334, w_035_014);
  or2  I044_120(w_044_120, w_033_012, w_024_025);
  not1 I044_127(w_044_127, w_000_114);
  and2 I044_130(w_044_130, w_016_046, w_021_061);
  not1 I044_133(w_044_133, w_026_328);
  or2  I044_136(w_044_136, w_024_069, w_011_284);
  or2  I044_140(w_044_140, w_005_216, w_039_113);
  nand2 I044_146(w_044_146, w_003_078, w_034_085);
  nand2 I044_151(w_044_151, w_042_040, w_029_154);
  or2  I044_153(w_044_153, w_015_088, w_015_040);
  nand2 I044_154(w_044_154, w_006_000, w_017_023);
  and2 I044_157(w_044_157, w_003_003, w_015_025);
  nand2 I044_158(w_044_158, w_020_012, w_037_078);
  and2 I044_161(w_044_161, w_019_036, w_031_000);
  not1 I044_163(w_044_163, w_010_291);
  nand2 I044_169(w_044_169, w_035_000, w_037_031);
  not1 I044_171(w_044_171, w_038_068);
  and2 I044_172(w_044_172, w_043_227, w_038_013);
  nand2 I044_184(w_044_184, w_014_241, w_030_148);
  not1 I044_193(w_044_193, w_024_176);
  nand2 I044_210(w_044_210, w_001_002, w_043_190);
  nand2 I044_212(w_044_212, w_024_295, w_027_232);
  nand2 I044_216(w_044_216, w_027_074, w_002_024);
  and2 I044_220(w_044_220, w_035_007, w_032_091);
  and2 I044_227(w_044_227, w_009_018, w_024_152);
  and2 I044_237(w_044_237, w_000_316, w_004_213);
  and2 I044_240(w_044_240, w_008_073, w_016_354);
  not1 I044_242(w_044_242, w_022_092);
  nand2 I044_245(w_044_245, w_006_000, w_016_354);
  not1 I044_258(w_044_258, w_018_155);
  nand2 I044_259(w_044_259, w_012_159, w_036_058);
  or2  I044_264(w_044_264, w_037_122, w_017_040);
  not1 I044_269(w_044_269, w_037_072);
  or2  I044_275(w_044_275, w_034_032, w_027_172);
  nand2 I044_277(w_044_277, w_026_294, w_015_113);
  and2 I044_281(w_044_281, w_002_006, w_009_131);
  nand2 I044_282(w_044_282, w_020_183, w_039_136);
  or2  I044_295(w_044_295, w_013_124, w_009_105);
  not1 I044_297(w_044_297, w_025_237);
  not1 I044_301(w_044_301, w_011_152);
  nand2 I044_302(w_044_302, w_025_240, w_005_090);
  and2 I044_307(w_044_307, w_042_193, w_022_071);
  or2  I044_323(w_044_323, w_003_006, w_039_346);
  not1 I044_326(w_044_326, w_007_125);
  or2  I045_001(w_045_001, w_027_400, w_017_093);
  not1 I045_004(w_045_004, w_041_125);
  or2  I045_005(w_045_005, w_027_354, w_017_037);
  not1 I045_008(w_045_008, w_018_297);
  nand2 I045_009(w_045_009, w_031_055, w_025_091);
  not1 I045_010(w_045_010, w_024_177);
  and2 I045_015(w_045_015, w_037_038, w_037_078);
  nand2 I045_018(w_045_018, w_035_083, w_007_095);
  nand2 I045_026(w_045_026, w_033_034, w_033_027);
  not1 I045_036(w_045_036, w_007_113);
  not1 I045_038(w_045_038, w_030_056);
  nand2 I045_039(w_045_039, w_016_053, w_008_283);
  not1 I045_065(w_045_065, w_003_003);
  and2 I045_066(w_045_066, w_012_041, w_029_130);
  or2  I045_069(w_045_069, w_028_232, w_020_042);
  or2  I045_082(w_045_082, w_024_121, w_015_085);
  and2 I045_090(w_045_090, w_044_038, w_025_093);
  or2  I045_092(w_045_092, w_016_020, w_031_020);
  not1 I045_094(w_045_094, w_015_083);
  nand2 I045_096(w_045_096, w_023_192, w_025_429);
  nand2 I045_099(w_045_099, w_001_001, w_027_070);
  not1 I045_103(w_045_103, w_007_183);
  or2  I045_104(w_045_104, w_018_096, w_037_067);
  and2 I045_106(w_045_106, w_009_161, w_003_076);
  or2  I045_112(w_045_112, w_030_085, w_039_400);
  nand2 I045_114(w_045_114, w_023_312, w_025_092);
  or2  I045_115(w_045_115, w_038_080, w_016_281);
  nand2 I045_118(w_045_118, w_006_000, w_023_233);
  not1 I045_119(w_045_119, w_013_097);
  not1 I045_125(w_045_125, w_026_127);
  not1 I045_132(w_045_132, w_042_102);
  and2 I045_135(w_045_135, w_003_005, w_033_007);
  not1 I045_136(w_045_136, w_029_019);
  nand2 I045_137(w_045_137, w_017_074, w_009_005);
  and2 I045_139(w_045_139, w_018_187, w_027_362);
  or2  I045_150(w_045_150, w_002_019, w_015_124);
  or2  I045_152(w_045_152, w_000_238, w_021_053);
  and2 I045_170(w_045_170, w_027_091, w_016_033);
  not1 I045_171(w_045_171, w_029_177);
  not1 I045_174(w_045_174, w_018_081);
  nand2 I045_177(w_045_177, w_037_001, w_041_129);
  nand2 I045_180(w_045_180, w_013_199, w_029_176);
  and2 I045_182(w_045_182, w_036_005, w_006_000);
  and2 I045_183(w_045_183, w_030_054, w_039_111);
  nand2 I045_184(w_045_184, w_003_025, w_035_032);
  nand2 I045_185(w_045_185, w_028_085, w_039_220);
  and2 I045_193(w_045_193, w_044_074, w_013_010);
  or2  I045_199(w_045_199, w_029_195, w_012_053);
  and2 I045_201(w_045_201, w_004_188, w_024_170);
  and2 I045_210(w_045_210, w_010_354, w_044_130);
  not1 I045_216(w_045_216, w_036_056);
  nand2 I045_229(w_045_229, w_023_285, w_034_170);
  not1 I045_231(w_045_231, w_005_185);
  or2  I045_241(w_045_241, w_002_002, w_015_131);
  nand2 I045_250(w_045_250, w_036_034, w_012_040);
  or2  I045_257(w_045_257, w_014_085, w_016_111);
  nand2 I045_276(w_045_276, w_009_228, w_027_114);
  and2 I045_283(w_045_283, w_044_140, w_001_000);
  and2 I045_284(w_045_284, w_030_196, w_008_270);
  and2 I046_004(w_046_004, w_001_002, w_018_322);
  nand2 I046_005(w_046_005, w_008_264, w_026_091);
  nand2 I046_006(w_046_006, w_010_020, w_001_005);
  and2 I046_007(w_046_007, w_014_236, w_026_072);
  or2  I046_008(w_046_008, w_038_002, w_019_043);
  or2  I046_010(w_046_010, w_004_032, w_037_140);
  not1 I046_011(w_046_011, w_032_072);
  and2 I046_015(w_046_015, w_003_054, w_004_017);
  nand2 I046_016(w_046_016, w_015_001, w_012_042);
  nand2 I046_021(w_046_021, w_043_212, w_033_048);
  or2  I046_023(w_046_023, w_000_328, w_003_019);
  nand2 I046_024(w_046_024, w_040_000, w_004_300);
  or2  I046_026(w_046_026, w_010_190, w_042_082);
  not1 I046_027(w_046_027, w_043_077);
  or2  I046_028(w_046_028, w_040_002, w_031_049);
  and2 I046_031(w_046_031, w_003_077, w_014_110);
  and2 I046_032(w_046_032, w_037_093, w_033_039);
  not1 I046_035(w_046_035, w_030_068);
  not1 I046_037(w_046_037, w_018_302);
  nand2 I046_039(w_046_039, w_028_017, w_034_043);
  nand2 I046_040(w_046_040, w_035_084, w_037_128);
  not1 I046_043(w_046_043, w_025_297);
  or2  I046_044(w_046_044, w_025_019, w_006_000);
  or2  I046_045(w_046_045, w_038_089, w_035_001);
  and2 I046_047(w_046_047, w_031_056, w_005_130);
  not1 I046_048(w_046_048, w_011_279);
  not1 I046_053(w_046_053, w_014_138);
  not1 I046_056(w_046_056, w_024_059);
  or2  I046_060(w_046_060, w_032_022, w_032_104);
  and2 I046_061(w_046_061, w_026_328, w_011_280);
  nand2 I046_062(w_046_062, w_021_003, w_038_089);
  not1 I046_063(w_046_063, w_017_143);
  not1 I046_067(w_046_067, w_019_015);
  not1 I046_084(w_046_084, w_006_000);
  and2 I046_086(w_046_086, w_025_264, w_001_003);
  nand2 I046_090(w_046_090, w_018_311, w_015_075);
  nand2 I046_094(w_046_094, w_022_081, w_008_072);
  or2  I046_097(w_046_097, w_021_030, w_019_029);
  and2 I046_107(w_046_107, w_035_108, w_008_048);
  not1 I046_108(w_046_108, w_020_012);
  and2 I046_113(w_046_113, w_041_141, w_012_256);
  not1 I046_114(w_046_114, w_041_175);
  and2 I046_115(w_046_115, w_016_005, w_032_171);
  and2 I046_118(w_046_118, w_001_004, w_039_046);
  and2 I046_119(w_046_119, w_019_020, w_005_088);
  not1 I046_122(w_046_122, w_045_174);
  and2 I046_125(w_046_125, w_028_370, w_042_170);
  or2  I046_126(w_046_126, w_000_250, w_021_101);
  or2  I046_127(w_046_127, w_043_237, w_039_463);
  nand2 I046_132(w_046_132, w_016_118, w_031_019);
  or2  I046_134(w_046_134, w_000_213, w_029_139);
  and2 I046_138(w_046_138, w_029_167, w_019_041);
  not1 I046_145(w_046_145, w_004_192);
  and2 I046_148(w_046_148, w_013_033, w_019_024);
  nand2 I046_150(w_046_150, w_004_474, w_039_100);
  not1 I046_151(w_046_151, w_026_018);
  or2  I046_161(w_046_161, w_024_178, w_025_071);
  not1 I046_165(w_046_165, w_045_066);
  nand2 I046_166(w_046_166, w_039_057, w_010_013);
  not1 I046_170(w_046_170, w_001_005);
  not1 I046_171(w_046_171, w_039_056);
  not1 I046_173(w_046_173, w_039_130);
  and2 I046_174(w_046_174, w_042_120, w_024_135);
  and2 I046_178(w_046_178, w_040_001, w_002_016);
  and2 I046_179(w_046_179, w_023_176, w_012_298);
  not1 I046_180(w_046_180, w_009_216);
  and2 I046_182(w_046_182, w_013_051, w_038_087);
  or2  I046_183(w_046_183, w_033_053, w_006_000);
  and2 I046_185(w_046_185, w_023_061, w_018_080);
  or2  I046_192(w_046_192, w_045_008, w_004_454);
  nand2 I046_198(w_046_198, w_040_000, w_039_357);
  and2 I046_208(w_046_208, w_002_010, w_023_050);
  nand2 I046_210(w_046_210, w_039_111, w_002_013);
  not1 I046_211(w_046_211, w_042_108);
  and2 I046_216(w_046_216, w_019_033, w_016_003);
  not1 I046_218(w_046_218, w_024_007);
  nand2 I046_221(w_046_221, w_027_005, w_024_008);
  not1 I047_001(w_047_001, w_007_128);
  nand2 I047_007(w_047_007, w_017_101, w_031_004);
  nand2 I047_013(w_047_013, w_001_006, w_043_226);
  and2 I047_015(w_047_015, w_028_076, w_037_047);
  not1 I047_022(w_047_022, w_002_018);
  nand2 I047_023(w_047_023, w_032_045, w_044_001);
  or2  I047_030(w_047_030, w_020_154, w_032_035);
  or2  I047_032(w_047_032, w_008_046, w_032_154);
  nand2 I047_036(w_047_036, w_017_177, w_005_094);
  nand2 I047_038(w_047_038, w_025_092, w_003_008);
  or2  I047_044(w_047_044, w_030_147, w_000_396);
  not1 I047_045(w_047_045, w_019_003);
  or2  I047_046(w_047_046, w_044_264, w_030_099);
  or2  I047_050(w_047_050, w_029_083, w_020_165);
  and2 I047_053(w_047_053, w_021_107, w_007_047);
  or2  I047_054(w_047_054, w_009_157, w_042_166);
  not1 I047_062(w_047_062, w_004_136);
  or2  I047_064(w_047_064, w_041_195, w_027_332);
  or2  I047_089(w_047_089, w_034_021, w_013_049);
  nand2 I047_090(w_047_090, w_009_067, w_032_025);
  and2 I047_102(w_047_102, w_003_059, w_002_001);
  not1 I047_103(w_047_103, w_017_177);
  nand2 I047_113(w_047_113, w_028_350, w_040_000);
  and2 I047_134(w_047_134, w_020_022, w_003_067);
  or2  I047_137(w_047_137, w_002_016, w_005_233);
  nand2 I047_141(w_047_141, w_011_131, w_013_151);
  not1 I047_151(w_047_151, w_014_113);
  and2 I047_152(w_047_152, w_032_030, w_036_105);
  nand2 I047_154(w_047_154, w_017_084, w_000_224);
  nand2 I047_162(w_047_162, w_022_005, w_011_336);
  and2 I047_164(w_047_164, w_003_065, w_002_019);
  nand2 I047_165(w_047_165, w_030_003, w_020_022);
  or2  I047_173(w_047_173, w_029_006, w_000_030);
  not1 I047_174(w_047_174, w_022_064);
  or2  I047_175(w_047_175, w_044_048, w_039_337);
  or2  I047_179(w_047_179, w_027_348, w_017_052);
  not1 I047_183(w_047_183, w_026_012);
  or2  I047_185(w_047_185, w_010_121, w_031_027);
  nand2 I047_196(w_047_196, w_033_008, w_005_071);
  or2  I047_201(w_047_201, w_046_127, w_029_083);
  not1 I047_202(w_047_202, w_038_030);
  not1 I047_207(w_047_207, w_032_077);
  or2  I047_216(w_047_216, w_003_076, w_036_046);
  nand2 I047_224(w_047_224, w_037_144, w_026_039);
  nand2 I047_228(w_047_228, w_031_050, w_032_034);
  not1 I047_229(w_047_229, w_001_002);
  or2  I047_230(w_047_230, w_043_222, w_035_001);
  or2  I047_231(w_047_231, w_040_000, w_014_198);
  and2 I047_233(w_047_233, w_019_005, w_013_047);
  and2 I047_234(w_047_234, w_017_179, w_041_235);
  or2  I047_235(w_047_235, w_005_017, w_018_054);
  nand2 I047_251(w_047_251, w_002_011, w_044_216);
  and2 I047_253(w_047_253, w_010_234, w_038_096);
  not1 I047_256(w_047_256, w_015_011);
  or2  I047_258(w_047_258, w_001_001, w_017_017);
  and2 I047_259(w_047_259, w_005_053, w_032_183);
  and2 I047_267(w_047_267, w_019_014, w_027_355);
  and2 I047_274(w_047_274, w_045_026, w_001_004);
  nand2 I047_276(w_047_276, w_012_278, w_009_016);
  nand2 I047_278(w_047_278, w_008_256, w_018_017);
  or2  I047_279(w_047_279, w_044_025, w_036_061);
  or2  I047_286(w_047_286, w_029_098, w_038_000);
  and2 I047_288(w_047_288, w_029_160, w_022_005);
  or2  I047_291(w_047_291, w_018_203, w_019_011);
  nand2 I047_292(w_047_292, w_027_404, w_004_003);
  not1 I047_293(w_047_293, w_021_106);
  and2 I047_306(w_047_306, w_039_331, w_019_029);
  or2  I047_310(w_047_310, w_039_117, w_038_041);
  not1 I047_316(w_047_316, w_035_029);
  nand2 I047_317(w_047_317, w_027_004, w_043_242);
  not1 I047_318(w_047_318, w_013_000);
  or2  I047_322(w_047_322, w_021_106, w_019_022);
  nand2 I047_329(w_047_329, w_031_037, w_020_066);
  and2 I047_330(w_047_330, w_043_179, w_038_046);
  nand2 I047_336(w_047_336, w_029_220, w_007_184);
  not1 I047_339(w_047_339, w_037_132);
  or2  I047_341(w_047_341, w_040_001, w_043_089);
  nand2 I047_350(w_047_350, w_004_310, w_042_047);
  nand2 I047_354(w_047_354, w_032_177, w_002_006);
  not1 I047_367(w_047_367, w_034_170);
  and2 I047_368(w_047_368, w_043_103, w_028_118);
  nand2 I047_390(w_047_390, w_045_185, w_046_171);
  and2 I047_397(w_047_397, w_025_195, w_035_015);
  and2 I047_400(w_047_400, w_003_016, w_005_203);
  nand2 I047_405(w_047_405, w_036_163, w_038_058);
  not1 I047_415(w_047_415, w_010_351);
  not1 I047_416(w_047_416, w_043_011);
  and2 I047_422(w_047_422, w_019_013, w_008_131);
  or2  I048_000(w_048_000, w_046_026, w_035_079);
  not1 I048_001(w_048_001, w_030_051);
  not1 I048_003(w_048_003, w_045_283);
  and2 I048_012(w_048_012, w_046_011, w_038_064);
  nand2 I048_014(w_048_014, w_028_386, w_034_093);
  and2 I048_019(w_048_019, w_017_016, w_046_063);
  and2 I048_020(w_048_020, w_037_090, w_042_188);
  nand2 I048_021(w_048_021, w_047_036, w_008_191);
  not1 I048_022(w_048_022, w_045_184);
  or2  I048_026(w_048_026, w_040_002, w_033_040);
  nand2 I048_029(w_048_029, w_019_045, w_038_066);
  and2 I048_033(w_048_033, w_021_034, w_033_046);
  nand2 I048_050(w_048_050, w_046_086, w_041_142);
  not1 I048_054(w_048_054, w_044_242);
  nand2 I048_055(w_048_055, w_017_144, w_042_223);
  not1 I048_056(w_048_056, w_011_169);
  and2 I048_061(w_048_061, w_016_130, w_020_115);
  nand2 I048_064(w_048_064, w_046_216, w_046_047);
  nand2 I048_071(w_048_071, w_020_186, w_025_101);
  nand2 I048_072(w_048_072, w_039_085, w_026_066);
  not1 I048_074(w_048_074, w_028_109);
  nand2 I048_079(w_048_079, w_038_077, w_033_020);
  or2  I048_081(w_048_081, w_033_010, w_005_161);
  and2 I048_083(w_048_083, w_010_260, w_045_250);
  and2 I048_085(w_048_085, w_023_284, w_042_005);
  and2 I048_087(w_048_087, w_016_175, w_021_029);
  nand2 I048_097(w_048_097, w_028_041, w_021_042);
  nand2 I048_100(w_048_100, w_005_026, w_034_085);
  not1 I048_103(w_048_103, w_039_216);
  not1 I048_104(w_048_104, w_028_334);
  not1 I048_107(w_048_107, w_008_311);
  nand2 I048_109(w_048_109, w_024_180, w_010_038);
  or2  I048_117(w_048_117, w_016_119, w_016_316);
  nand2 I048_118(w_048_118, w_026_034, w_019_022);
  not1 I048_119(w_048_119, w_018_137);
  not1 I048_128(w_048_128, w_015_015);
  not1 I048_132(w_048_132, w_011_031);
  and2 I048_133(w_048_133, w_036_120, w_002_003);
  nand2 I048_137(w_048_137, w_037_125, w_006_000);
  nand2 I048_143(w_048_143, w_013_239, w_025_456);
  nand2 I048_147(w_048_147, w_002_022, w_033_024);
  nand2 I048_149(w_048_149, w_025_249, w_043_121);
  or2  I048_169(w_048_169, w_015_070, w_001_002);
  not1 I048_171(w_048_171, w_009_154);
  not1 I048_184(w_048_184, w_018_135);
  nand2 I048_187(w_048_187, w_012_012, w_031_040);
  not1 I048_190(w_048_190, w_014_025);
  not1 I048_193(w_048_193, w_034_124);
  nand2 I048_196(w_048_196, w_017_051, w_037_089);
  nand2 I048_207(w_048_207, w_021_010, w_026_113);
  and2 I048_209(w_048_209, w_024_110, w_036_200);
  nand2 I048_211(w_048_211, w_030_138, w_015_095);
  nand2 I048_216(w_048_216, w_012_074, w_043_099);
  or2  I048_233(w_048_233, w_014_110, w_030_098);
  not1 I048_234(w_048_234, w_029_116);
  and2 I048_247(w_048_247, w_002_001, w_042_094);
  nand2 I048_255(w_048_255, w_044_193, w_038_019);
  or2  I048_265(w_048_265, w_018_089, w_003_091);
  and2 I048_268(w_048_268, w_017_085, w_017_111);
  or2  I048_271(w_048_271, w_006_000, w_038_032);
  or2  I048_279(w_048_279, w_047_183, w_005_094);
  nand2 I048_280(w_048_280, w_017_141, w_021_023);
  or2  I048_281(w_048_281, w_024_185, w_014_104);
  and2 I048_284(w_048_284, w_014_134, w_009_018);
  nand2 I048_285(w_048_285, w_042_265, w_038_081);
  nand2 I048_303(w_048_303, w_012_161, w_033_054);
  nand2 I048_304(w_048_304, w_043_183, w_001_004);
  or2  I048_314(w_048_314, w_009_032, w_004_080);
  and2 I048_317(w_048_317, w_047_276, w_005_127);
  nand2 I048_342(w_048_342, w_020_050, w_015_116);
  and2 I048_347(w_048_347, w_027_449, w_026_151);
  or2  I048_355(w_048_355, w_006_000, w_021_028);
  not1 I048_366(w_048_366, w_029_128);
  nand2 I049_000(w_049_000, w_002_000, w_021_060);
  not1 I049_002(w_049_002, w_019_022);
  not1 I049_003(w_049_003, w_030_135);
  or2  I049_008(w_049_008, w_033_009, w_043_080);
  nand2 I049_012(w_049_012, w_043_192, w_007_171);
  or2  I049_023(w_049_023, w_039_306, w_016_038);
  not1 I049_025(w_049_025, w_006_000);
  and2 I049_030(w_049_030, w_006_000, w_018_124);
  nand2 I049_038(w_049_038, w_042_160, w_033_040);
  not1 I049_044(w_049_044, w_038_056);
  or2  I049_047(w_049_047, w_015_005, w_003_080);
  and2 I049_060(w_049_060, w_038_040, w_038_001);
  and2 I049_065(w_049_065, w_020_163, w_021_024);
  or2  I049_066(w_049_066, w_015_034, w_005_093);
  and2 I049_070(w_049_070, w_037_015, w_047_179);
  and2 I049_071(w_049_071, w_002_001, w_048_087);
  nand2 I049_074(w_049_074, w_020_152, w_007_175);
  and2 I049_076(w_049_076, w_046_048, w_035_090);
  or2  I049_079(w_049_079, w_039_496, w_027_154);
  or2  I049_087(w_049_087, w_047_291, w_037_066);
  and2 I049_090(w_049_090, w_021_034, w_040_002);
  and2 I049_091(w_049_091, w_006_000, w_011_197);
  or2  I049_100(w_049_100, w_046_174, w_007_371);
  not1 I049_107(w_049_107, w_032_085);
  not1 I049_108(w_049_108, w_009_032);
  and2 I049_113(w_049_113, w_000_132, w_034_182);
  nand2 I049_121(w_049_121, w_016_185, w_011_327);
  not1 I049_137(w_049_137, w_028_255);
  or2  I049_139(w_049_139, w_029_234, w_021_057);
  not1 I049_149(w_049_149, w_029_075);
  and2 I049_165(w_049_165, w_042_002, w_008_063);
  not1 I049_166(w_049_166, w_017_054);
  nand2 I049_173(w_049_173, w_018_050, w_015_060);
  or2  I049_174(w_049_174, w_020_094, w_011_031);
  not1 I049_179(w_049_179, w_009_040);
  not1 I049_182(w_049_182, w_041_003);
  not1 I049_185(w_049_185, w_035_018);
  nand2 I049_189(w_049_189, w_027_020, w_003_099);
  not1 I049_191(w_049_191, w_013_122);
  or2  I049_200(w_049_200, w_046_179, w_017_146);
  nand2 I049_201(w_049_201, w_004_019, w_019_049);
  not1 I049_218(w_049_218, w_006_000);
  or2  I049_219(w_049_219, w_037_124, w_041_011);
  and2 I049_231(w_049_231, w_039_001, w_014_229);
  and2 I049_244(w_049_244, w_014_206, w_027_347);
  or2  I049_250(w_049_250, w_007_177, w_046_037);
  nand2 I049_262(w_049_262, w_028_360, w_008_274);
  and2 I049_266(w_049_266, w_022_148, w_026_197);
  and2 I049_272(w_049_272, w_032_069, w_021_100);
  and2 I049_273(w_049_273, w_048_149, w_002_004);
  nand2 I049_277(w_049_277, w_002_006, w_018_045);
  and2 I049_285(w_049_285, w_019_005, w_005_012);
  and2 I049_297(w_049_297, w_047_054, w_002_026);
  or2  I049_301(w_049_301, w_040_001, w_041_169);
  and2 I049_307(w_049_307, w_031_044, w_004_080);
  not1 I049_320(w_049_320, w_026_042);
  or2  I049_323(w_049_323, w_007_404, w_047_339);
  not1 I049_329(w_049_329, w_007_159);
  not1 I049_333(w_049_333, w_042_221);
  not1 I049_338(w_049_338, w_034_061);
  nand2 I049_343(w_049_343, w_014_073, w_002_008);
  or2  I049_347(w_049_347, w_045_132, w_029_182);
  not1 I049_361(w_049_361, w_035_040);
  and2 I049_377(w_049_377, w_003_044, w_027_135);
  and2 I049_380(w_049_380, w_028_056, w_008_090);
  nand2 I049_383(w_049_383, w_038_062, w_007_030);
  nand2 I049_388(w_049_388, w_045_103, w_038_044);
  nand2 I049_400(w_049_400, w_018_142, w_024_088);
  and2 I049_401(w_049_401, w_038_044, w_021_106);
  and2 I049_403(w_049_403, w_008_043, w_038_035);
  and2 I050_001(w_050_001, w_034_088, w_013_099);
  nand2 I050_002(w_050_002, w_005_021, w_003_085);
  or2  I050_003(w_050_003, w_025_362, w_018_132);
  and2 I050_007(w_050_007, w_023_373, w_012_026);
  nand2 I050_008(w_050_008, w_026_361, w_031_007);
  nand2 I050_009(w_050_009, w_036_272, w_038_008);
  not1 I050_010(w_050_010, w_006_000);
  or2  I050_014(w_050_014, w_040_006, w_020_031);
  and2 I050_015(w_050_015, w_003_053, w_005_239);
  not1 I050_016(w_050_016, w_043_202);
  and2 I050_017(w_050_017, w_002_017, w_032_034);
  or2  I050_022(w_050_022, w_007_069, w_047_102);
  nand2 I050_026(w_050_026, w_038_070, w_011_100);
  not1 I050_030(w_050_030, w_010_041);
  or2  I050_034(w_050_034, w_019_017, w_024_188);
  nand2 I050_035(w_050_035, w_046_084, w_040_001);
  or2  I050_038(w_050_038, w_048_026, w_014_002);
  nand2 I050_039(w_050_039, w_026_276, w_026_302);
  not1 I050_042(w_050_042, w_022_044);
  and2 I050_043(w_050_043, w_014_092, w_024_124);
  nand2 I050_045(w_050_045, w_014_184, w_027_232);
  nand2 I050_046(w_050_046, w_005_008, w_045_257);
  nand2 I050_047(w_050_047, w_048_133, w_040_006);
  not1 I050_051(w_050_051, w_024_021);
  not1 I050_052(w_050_052, w_003_049);
  and2 I050_054(w_050_054, w_009_063, w_044_032);
  and2 I050_055(w_050_055, w_013_149, w_034_254);
  and2 I050_057(w_050_057, w_046_192, w_033_039);
  nand2 I050_058(w_050_058, w_040_000, w_027_007);
  nand2 I050_060(w_050_060, w_023_210, w_032_188);
  not1 I050_063(w_050_063, w_005_080);
  and2 I050_067(w_050_067, w_011_098, w_007_066);
  nand2 I050_070(w_050_070, w_043_000, w_016_019);
  nand2 I050_073(w_050_073, w_022_020, w_034_200);
  and2 I050_087(w_050_087, w_026_162, w_011_052);
  or2  I050_096(w_050_096, w_027_185, w_049_401);
  or2  I050_102(w_050_102, w_031_042, w_012_027);
  and2 I050_106(w_050_106, w_018_285, w_041_139);
  not1 I050_111(w_050_111, w_040_005);
  or2  I050_112(w_050_112, w_031_030, w_014_150);
  nand2 I050_113(w_050_113, w_007_141, w_002_008);
  and2 I050_117(w_050_117, w_014_091, w_011_159);
  and2 I050_121(w_050_121, w_016_176, w_026_088);
  and2 I050_124(w_050_124, w_042_275, w_037_120);
  or2  I050_125(w_050_125, w_020_159, w_000_287);
  or2  I050_126(w_050_126, w_035_056, w_040_000);
  nand2 I050_128(w_050_128, w_013_108, w_039_145);
  and2 I050_136(w_050_136, w_015_040, w_040_005);
  and2 I050_138(w_050_138, w_024_068, w_012_109);
  and2 I050_142(w_050_142, w_031_036, w_022_021);
  not1 I050_146(w_050_146, w_019_007);
  or2  I050_149(w_050_149, w_048_097, w_049_121);
  and2 I050_152(w_050_152, w_022_127, w_049_400);
  or2  I050_155(w_050_155, w_044_212, w_008_315);
  and2 I050_161(w_050_161, w_015_006, w_033_003);
  or2  I050_172(w_050_172, w_042_051, w_005_177);
  not1 I050_173(w_050_173, w_026_038);
  or2  I050_174(w_050_174, w_042_075, w_034_008);
  or2  I050_175(w_050_175, w_014_234, w_024_089);
  or2  I050_176(w_050_176, w_033_000, w_008_154);
  or2  I050_180(w_050_180, w_041_031, w_018_183);
  and2 I050_182(w_050_182, w_031_036, w_043_211);
  and2 I050_184(w_050_184, w_003_086, w_028_074);
  and2 I050_187(w_050_187, w_035_090, w_006_000);
  or2  I050_188(w_050_188, w_012_005, w_019_043);
  nand2 I050_192(w_050_192, w_035_007, w_027_239);
  not1 I050_193(w_050_193, w_045_136);
  nand2 I050_198(w_050_198, w_049_377, w_003_012);
  and2 I050_199(w_050_199, w_040_003, w_026_131);
  and2 I050_204(w_050_204, w_026_099, w_030_026);
  or2  I051_001(w_051_001, w_018_119, w_012_277);
  or2  I051_002(w_051_002, w_007_168, w_043_101);
  and2 I051_003(w_051_003, w_007_104, w_010_191);
  or2  I051_008(w_051_008, w_008_209, w_024_235);
  nand2 I051_010(w_051_010, w_015_004, w_021_015);
  and2 I051_016(w_051_016, w_000_014, w_037_022);
  not1 I051_017(w_051_017, w_033_051);
  not1 I051_018(w_051_018, w_007_101);
  and2 I051_023(w_051_023, w_005_014, w_011_117);
  not1 I051_026(w_051_026, w_038_051);
  nand2 I051_028(w_051_028, w_048_169, w_012_126);
  not1 I051_031(w_051_031, w_010_027);
  not1 I051_033(w_051_033, w_010_015);
  or2  I051_035(w_051_035, w_043_156, w_049_074);
  or2  I051_041(w_051_041, w_012_132, w_020_172);
  or2  I051_042(w_051_042, w_019_001, w_020_037);
  and2 I051_045(w_051_045, w_026_227, w_004_021);
  not1 I051_046(w_051_046, w_033_042);
  and2 I051_056(w_051_056, w_017_074, w_022_101);
  and2 I051_060(w_051_060, w_029_237, w_010_276);
  and2 I051_076(w_051_076, w_030_191, w_040_004);
  or2  I051_078(w_051_078, w_014_166, w_035_011);
  and2 I051_081(w_051_081, w_046_094, w_030_085);
  and2 I051_085(w_051_085, w_047_053, w_022_034);
  or2  I051_094(w_051_094, w_044_158, w_038_047);
  and2 I051_095(w_051_095, w_007_146, w_037_013);
  or2  I051_097(w_051_097, w_013_110, w_040_000);
  nand2 I051_098(w_051_098, w_034_108, w_032_145);
  not1 I051_101(w_051_101, w_045_135);
  nand2 I051_104(w_051_104, w_001_003, w_010_201);
  or2  I051_107(w_051_107, w_047_103, w_031_032);
  not1 I051_110(w_051_110, w_025_336);
  or2  I051_117(w_051_117, w_042_202, w_007_215);
  nand2 I051_119(w_051_119, w_046_165, w_050_009);
  nand2 I051_124(w_051_124, w_003_057, w_005_181);
  not1 I051_128(w_051_128, w_013_066);
  and2 I051_130(w_051_130, w_049_087, w_031_003);
  or2  I051_132(w_051_132, w_008_023, w_018_259);
  nand2 I051_146(w_051_146, w_000_014, w_044_053);
  and2 I051_151(w_051_151, w_030_010, w_018_246);
  not1 I051_153(w_051_153, w_007_248);
  not1 I051_154(w_051_154, w_025_445);
  or2  I051_159(w_051_159, w_034_271, w_035_078);
  not1 I051_164(w_051_164, w_029_063);
  not1 I051_165(w_051_165, w_016_011);
  not1 I051_172(w_051_172, w_012_077);
  not1 I051_181(w_051_181, w_005_238);
  and2 I051_182(w_051_182, w_047_310, w_032_018);
  and2 I051_197(w_051_197, w_031_037, w_003_079);
  not1 I051_198(w_051_198, w_040_000);
  and2 I051_210(w_051_210, w_028_029, w_038_077);
  or2  I051_211(w_051_211, w_034_093, w_025_375);
  or2  I051_218(w_051_218, w_038_079, w_000_122);
  or2  I051_221(w_051_221, w_040_001, w_039_348);
  and2 I051_223(w_051_223, w_040_003, w_012_249);
  not1 I051_226(w_051_226, w_030_081);
  or2  I051_238(w_051_238, w_014_181, w_040_002);
  nand2 I051_246(w_051_246, w_004_462, w_004_191);
  not1 I051_253(w_051_253, w_007_124);
  nand2 I051_260(w_051_260, w_047_007, w_047_230);
  or2  I051_266(w_051_266, w_028_284, w_001_006);
  or2  I051_286(w_051_286, w_038_023, w_037_118);
  nand2 I051_306(w_051_306, w_011_056, w_011_287);
  nand2 I051_313(w_051_313, w_048_268, w_016_349);
  nand2 I052_004(w_052_004, w_035_002, w_037_059);
  or2  I052_005(w_052_005, w_017_098, w_016_356);
  nand2 I052_006(w_052_006, w_004_021, w_000_158);
  nand2 I052_007(w_052_007, w_011_224, w_051_153);
  not1 I052_008(w_052_008, w_048_255);
  or2  I052_009(w_052_009, w_046_113, w_034_100);
  or2  I052_012(w_052_012, w_023_002, w_046_198);
  and2 I052_013(w_052_013, w_026_048, w_044_154);
  nand2 I052_015(w_052_015, w_037_091, w_044_109);
  or2  I052_016(w_052_016, w_027_325, w_011_001);
  and2 I052_017(w_052_017, w_004_111, w_012_034);
  or2  I052_018(w_052_018, w_014_245, w_034_042);
  or2  I052_019(w_052_019, w_027_154, w_011_095);
  nand2 I052_020(w_052_020, w_000_259, w_036_184);
  or2  I052_022(w_052_022, w_020_014, w_042_255);
  and2 I052_023(w_052_023, w_014_227, w_039_435);
  nand2 I052_027(w_052_027, w_014_193, w_009_103);
  and2 I052_033(w_052_033, w_026_248, w_024_196);
  not1 I052_034(w_052_034, w_009_037);
  nand2 I052_035(w_052_035, w_003_090, w_002_019);
  not1 I052_036(w_052_036, w_014_140);
  nand2 I052_038(w_052_038, w_039_381, w_007_049);
  or2  I052_039(w_052_039, w_019_025, w_023_013);
  and2 I052_040(w_052_040, w_049_113, w_020_037);
  or2  I052_047(w_052_047, w_037_115, w_034_179);
  or2  I052_048(w_052_048, w_019_018, w_014_083);
  or2  I052_049(w_052_049, w_022_095, w_010_241);
  not1 I052_051(w_052_051, w_022_123);
  nand2 I052_054(w_052_054, w_051_085, w_001_005);
  and2 I052_056(w_052_056, w_037_052, w_030_022);
  nand2 I052_058(w_052_058, w_041_241, w_049_361);
  not1 I052_061(w_052_061, w_047_038);
  nand2 I052_066(w_052_066, w_037_064, w_033_052);
  nand2 I052_068(w_052_068, w_030_080, w_035_065);
  or2  I052_071(w_052_071, w_044_237, w_035_017);
  not1 I052_084(w_052_084, w_017_012);
  not1 I052_085(w_052_085, w_040_006);
  nand2 I052_086(w_052_086, w_043_094, w_040_003);
  not1 I052_095(w_052_095, w_027_235);
  and2 I052_097(w_052_097, w_014_119, w_027_010);
  or2  I052_098(w_052_098, w_047_046, w_050_010);
  and2 I052_101(w_052_101, w_025_190, w_038_010);
  nand2 I052_103(w_052_103, w_012_374, w_022_069);
  nand2 I052_104(w_052_104, w_044_014, w_049_262);
  and2 I052_110(w_052_110, w_009_090, w_015_113);
  nand2 I052_112(w_052_112, w_023_122, w_003_034);
  not1 I052_113(w_052_113, w_005_244);
  and2 I052_115(w_052_115, w_030_077, w_012_073);
  or2  I052_116(w_052_116, w_015_122, w_031_054);
  or2  I053_000(w_053_000, w_016_260, w_003_003);
  not1 I053_001(w_053_001, w_016_297);
  and2 I053_002(w_053_002, w_039_295, w_049_091);
  and2 I053_003(w_053_003, w_047_233, w_050_198);
  or2  I053_004(w_053_004, w_051_182, w_034_194);
  and2 I053_005(w_053_005, w_041_147, w_013_155);
  and2 I053_006(w_053_006, w_046_056, w_045_092);
  not1 I053_007(w_053_007, w_048_355);
  nand2 I053_009(w_053_009, w_006_000, w_028_215);
  nand2 I053_011(w_053_011, w_002_020, w_046_185);
  nand2 I053_013(w_053_013, w_035_069, w_018_212);
  not1 I053_014(w_053_014, w_046_067);
  nand2 I053_015(w_053_015, w_016_071, w_048_100);
  nand2 I053_016(w_053_016, w_033_058, w_005_158);
  or2  I053_018(w_053_018, w_011_249, w_018_022);
  and2 I053_019(w_053_019, w_007_022, w_049_285);
  and2 I053_021(w_053_021, w_004_272, w_020_001);
  or2  I053_022(w_053_022, w_050_180, w_040_001);
  and2 I053_023(w_053_023, w_047_291, w_009_121);
  nand2 I053_025(w_053_025, w_023_014, w_043_056);
  and2 I053_026(w_053_026, w_050_016, w_027_203);
  not1 I053_027(w_053_027, w_018_235);
  nand2 I053_028(w_053_028, w_017_083, w_042_178);
  and2 I053_029(w_053_029, w_008_131, w_024_251);
  nand2 I053_031(w_053_031, w_042_072, w_008_047);
  not1 I053_033(w_053_033, w_022_096);
  nand2 I053_034(w_053_034, w_016_349, w_039_002);
  and2 I053_035(w_053_035, w_003_027, w_036_008);
  nand2 I053_037(w_053_037, w_025_265, w_016_315);
  not1 I053_039(w_053_039, w_037_002);
  and2 I054_000(w_054_000, w_002_011, w_029_024);
  and2 I054_003(w_054_003, w_024_185, w_002_000);
  not1 I054_005(w_054_005, w_006_000);
  and2 I054_012(w_054_012, w_006_000, w_034_278);
  nand2 I054_013(w_054_013, w_041_150, w_047_317);
  nand2 I054_014(w_054_014, w_008_046, w_013_148);
  and2 I054_015(w_054_015, w_006_000, w_046_016);
  nand2 I054_018(w_054_018, w_023_379, w_000_189);
  or2  I054_020(w_054_020, w_015_027, w_035_009);
  and2 I054_023(w_054_023, w_038_020, w_022_014);
  nand2 I054_029(w_054_029, w_009_012, w_006_000);
  or2  I054_030(w_054_030, w_003_100, w_003_072);
  and2 I054_031(w_054_031, w_018_297, w_005_121);
  or2  I054_034(w_054_034, w_005_052, w_036_205);
  not1 I054_038(w_054_038, w_018_015);
  not1 I054_040(w_054_040, w_008_077);
  nand2 I054_042(w_054_042, w_050_096, w_028_254);
  or2  I054_043(w_054_043, w_031_017, w_024_173);
  or2  I054_044(w_054_044, w_038_024, w_016_362);
  or2  I054_048(w_054_048, w_017_166, w_053_007);
  nand2 I054_051(w_054_051, w_025_416, w_038_064);
  or2  I054_054(w_054_054, w_042_134, w_050_125);
  and2 I054_055(w_054_055, w_016_391, w_018_026);
  nand2 I054_056(w_054_056, w_007_333, w_049_333);
  nand2 I054_057(w_054_057, w_038_008, w_047_062);
  nand2 I054_063(w_054_063, w_011_230, w_027_128);
  or2  I054_064(w_054_064, w_014_252, w_017_049);
  nand2 I054_068(w_054_068, w_039_344, w_010_144);
  not1 I054_070(w_054_070, w_048_107);
  and2 I054_073(w_054_073, w_040_003, w_002_006);
  or2  I054_074(w_054_074, w_049_277, w_007_174);
  or2  I054_081(w_054_081, w_051_098, w_040_003);
  not1 I054_083(w_054_083, w_013_172);
  not1 I054_084(w_054_084, w_015_096);
  or2  I054_088(w_054_088, w_050_054, w_022_072);
  not1 I054_089(w_054_089, w_019_034);
  nand2 I054_090(w_054_090, w_032_171, w_044_094);
  or2  I054_097(w_054_097, w_030_076, w_029_153);
  and2 I054_100(w_054_100, w_007_382, w_042_152);
  not1 I054_101(w_054_101, w_047_306);
  not1 I054_106(w_054_106, w_042_113);
  and2 I054_110(w_054_110, w_013_061, w_005_135);
  not1 I054_113(w_054_113, w_017_047);
  nand2 I054_115(w_054_115, w_015_037, w_041_295);
  and2 I054_118(w_054_118, w_049_044, w_018_095);
  not1 I054_125(w_054_125, w_022_114);
  or2  I054_134(w_054_134, w_011_194, w_019_004);
  and2 I054_137(w_054_137, w_046_031, w_018_059);
  and2 I054_146(w_054_146, w_047_001, w_035_028);
  not1 I054_165(w_054_165, w_004_356);
  not1 I054_166(w_054_166, w_041_048);
  nand2 I054_170(w_054_170, w_015_027, w_038_094);
  and2 I054_172(w_054_172, w_030_189, w_028_323);
  or2  I054_177(w_054_177, w_032_143, w_029_173);
  or2  I054_178(w_054_178, w_014_204, w_039_496);
  or2  I054_191(w_054_191, w_035_008, w_016_294);
  and2 I054_199(w_054_199, w_019_033, w_001_002);
  not1 I054_204(w_054_204, w_016_336);
  or2  I054_205(w_054_205, w_037_089, w_046_097);
  nand2 I054_208(w_054_208, w_038_099, w_048_255);
  nand2 I054_210(w_054_210, w_024_196, w_043_065);
  not1 I054_211(w_054_211, w_021_042);
  nand2 I055_000(w_055_000, w_013_229, w_054_137);
  or2  I055_001(w_055_001, w_028_237, w_033_029);
  or2  I055_002(w_055_002, w_046_005, w_044_032);
  not1 I055_005(w_055_005, w_017_027);
  nand2 I055_011(w_055_011, w_023_244, w_003_073);
  or2  I055_012(w_055_012, w_045_010, w_016_044);
  nand2 I055_016(w_055_016, w_005_065, w_007_347);
  and2 I055_018(w_055_018, w_053_037, w_024_111);
  or2  I055_019(w_055_019, w_049_023, w_024_009);
  not1 I055_022(w_055_022, w_039_397);
  not1 I055_028(w_055_028, w_047_229);
  not1 I055_029(w_055_029, w_038_016);
  and2 I055_031(w_055_031, w_032_055, w_020_096);
  nand2 I055_033(w_055_033, w_050_060, w_044_037);
  nand2 I055_035(w_055_035, w_022_067, w_007_347);
  nand2 I055_036(w_055_036, w_042_096, w_005_167);
  not1 I055_037(w_055_037, w_035_018);
  nand2 I055_039(w_055_039, w_012_248, w_035_045);
  nand2 I055_040(w_055_040, w_017_027, w_028_308);
  and2 I055_043(w_055_043, w_039_268, w_011_319);
  and2 I055_045(w_055_045, w_021_067, w_004_393);
  nand2 I055_046(w_055_046, w_039_404, w_016_223);
  and2 I055_047(w_055_047, w_031_043, w_048_187);
  and2 I055_048(w_055_048, w_044_028, w_029_052);
  and2 I055_049(w_055_049, w_040_006, w_014_133);
  and2 I055_051(w_055_051, w_011_232, w_043_060);
  or2  I055_052(w_055_052, w_020_159, w_007_118);
  or2  I055_053(w_055_053, w_008_154, w_052_015);
  or2  I055_055(w_055_055, w_042_131, w_032_002);
  or2  I055_056(w_055_056, w_025_376, w_046_061);
  nand2 I055_059(w_055_059, w_053_029, w_022_064);
  or2  I055_064(w_055_064, w_014_028, w_014_174);
  nand2 I055_065(w_055_065, w_038_014, w_052_006);
  or2  I055_068(w_055_068, w_007_116, w_021_039);
  nand2 I055_069(w_055_069, w_023_071, w_039_104);
  and2 I055_071(w_055_071, w_016_285, w_004_308);
  or2  I055_072(w_055_072, w_032_096, w_029_044);
  or2  I055_074(w_055_074, w_003_032, w_034_170);
  not1 I055_075(w_055_075, w_000_173);
  not1 I055_076(w_055_076, w_024_244);
  and2 I055_077(w_055_077, w_015_049, w_000_391);
  or2  I055_078(w_055_078, w_017_059, w_038_073);
  or2  I055_079(w_055_079, w_039_338, w_006_000);
  and2 I055_083(w_055_083, w_013_189, w_025_331);
  or2  I055_085(w_055_085, w_002_020, w_036_163);
  not1 I055_086(w_055_086, w_042_088);
  or2  I056_003(w_056_003, w_046_053, w_029_040);
  nand2 I056_008(w_056_008, w_038_070, w_021_033);
  nand2 I056_010(w_056_010, w_029_095, w_024_073);
  and2 I056_015(w_056_015, w_030_090, w_055_033);
  not1 I056_020(w_056_020, w_052_113);
  not1 I056_026(w_056_026, w_032_110);
  nand2 I056_036(w_056_036, w_016_002, w_001_001);
  or2  I056_043(w_056_043, w_049_000, w_055_075);
  nand2 I056_046(w_056_046, w_023_231, w_048_281);
  not1 I056_047(w_056_047, w_024_164);
  not1 I056_048(w_056_048, w_055_036);
  and2 I056_050(w_056_050, w_022_004, w_045_241);
  nand2 I056_053(w_056_053, w_048_314, w_003_093);
  or2  I056_054(w_056_054, w_027_115, w_023_238);
  nand2 I056_056(w_056_056, w_007_087, w_051_035);
  nand2 I056_058(w_056_058, w_028_382, w_014_014);
  or2  I056_063(w_056_063, w_039_395, w_047_064);
  nand2 I056_068(w_056_068, w_047_341, w_029_047);
  not1 I056_071(w_056_071, w_031_010);
  not1 I056_074(w_056_074, w_035_002);
  and2 I056_076(w_056_076, w_000_353, w_023_402);
  not1 I056_078(w_056_078, w_022_112);
  nand2 I056_087(w_056_087, w_009_177, w_035_039);
  or2  I056_092(w_056_092, w_046_008, w_025_214);
  and2 I056_093(w_056_093, w_007_035, w_035_107);
  and2 I056_100(w_056_100, w_030_101, w_034_084);
  or2  I056_102(w_056_102, w_005_153, w_023_386);
  or2  I056_105(w_056_105, w_003_052, w_047_397);
  and2 I056_106(w_056_106, w_027_063, w_053_035);
  nand2 I056_109(w_056_109, w_016_263, w_043_121);
  not1 I056_110(w_056_110, w_044_007);
  or2  I056_111(w_056_111, w_017_058, w_054_170);
  nand2 I056_118(w_056_118, w_029_179, w_021_052);
  nand2 I056_121(w_056_121, w_006_000, w_017_133);
  or2  I056_122(w_056_122, w_022_016, w_016_173);
  or2  I056_131(w_056_131, w_039_067, w_004_315);
  nand2 I056_137(w_056_137, w_014_063, w_044_240);
  nand2 I056_138(w_056_138, w_040_002, w_026_283);
  or2  I056_139(w_056_139, w_041_155, w_034_240);
  or2  I056_141(w_056_141, w_012_014, w_043_016);
  and2 I056_142(w_056_142, w_026_035, w_034_223);
  and2 I056_143(w_056_143, w_029_161, w_039_274);
  and2 I056_146(w_056_146, w_027_427, w_019_020);
  not1 I056_147(w_056_147, w_045_094);
  nand2 I056_148(w_056_148, w_001_003, w_042_158);
  or2  I056_149(w_056_149, w_012_336, w_047_152);
  nand2 I056_151(w_056_151, w_038_040, w_011_140);
  nand2 I056_162(w_056_162, w_008_125, w_001_003);
  and2 I056_163(w_056_163, w_050_111, w_020_175);
  and2 I056_164(w_056_164, w_031_061, w_012_300);
  nand2 I056_169(w_056_169, w_033_001, w_036_095);
  not1 I056_170(w_056_170, w_040_001);
  or2  I056_175(w_056_175, w_013_014, w_010_345);
  nand2 I056_176(w_056_176, w_030_093, w_020_056);
  nand2 I056_177(w_056_177, w_034_262, w_010_023);
  or2  I057_001(w_057_001, w_017_008, w_011_123);
  nand2 I057_002(w_057_002, w_040_003, w_009_079);
  not1 I057_003(w_057_003, w_036_168);
  not1 I057_004(w_057_004, w_035_079);
  or2  I057_005(w_057_005, w_008_018, w_050_149);
  or2  I057_006(w_057_006, w_031_037, w_049_231);
  or2  I057_007(w_057_007, w_033_033, w_047_390);
  nand2 I057_008(w_057_008, w_007_250, w_014_116);
  not1 I057_010(w_057_010, w_056_121);
  and2 I057_011(w_057_011, w_034_122, w_007_072);
  or2  I057_012(w_057_012, w_017_073, w_038_011);
  or2  I057_015(w_057_015, w_027_009, w_002_005);
  or2  I057_016(w_057_016, w_056_175, w_025_446);
  and2 I057_018(w_057_018, w_048_119, w_007_026);
  and2 I057_019(w_057_019, w_004_198, w_031_032);
  not1 I057_020(w_057_020, w_003_003);
  nand2 I057_021(w_057_021, w_023_272, w_002_021);
  and2 I057_022(w_057_022, w_004_110, w_035_057);
  and2 I057_023(w_057_023, w_003_015, w_033_035);
  not1 I057_024(w_057_024, w_017_052);
  not1 I057_027(w_057_027, w_050_199);
  and2 I057_028(w_057_028, w_041_207, w_029_095);
  and2 I057_030(w_057_030, w_053_028, w_006_000);
  or2  I057_031(w_057_031, w_049_383, w_032_039);
  not1 I057_033(w_057_033, w_024_051);
  and2 I057_034(w_057_034, w_017_071, w_050_008);
  nand2 I057_035(w_057_035, w_039_160, w_052_110);
  nand2 I057_036(w_057_036, w_044_184, w_034_145);
  not1 I057_037(w_057_037, w_040_002);
  and2 I057_039(w_057_039, w_056_146, w_027_256);
  not1 I057_041(w_057_041, w_012_263);
  or2  I057_044(w_057_044, w_026_013, w_017_171);
  and2 I057_046(w_057_046, w_028_052, w_005_097);
  nand2 I057_048(w_057_048, w_007_186, w_022_076);
  and2 I057_049(w_057_049, w_052_017, w_039_370);
  nand2 I057_050(w_057_050, w_021_089, w_027_186);
  nand2 I057_051(w_057_051, w_044_049, w_051_181);
  and2 I057_052(w_057_052, w_036_201, w_038_012);
  nand2 I057_053(w_057_053, w_030_086, w_018_075);
  not1 I057_054(w_057_054, w_013_050);
  nand2 I057_056(w_057_056, w_034_067, w_031_040);
  nand2 I057_057(w_057_057, w_017_159, w_012_083);
  and2 I057_058(w_057_058, w_023_050, w_011_282);
  nand2 I057_059(w_057_059, w_008_058, w_044_157);
  and2 I057_060(w_057_060, w_022_084, w_015_051);
  not1 I058_000(w_058_000, w_051_128);
  not1 I058_001(w_058_001, w_034_139);
  nand2 I058_005(w_058_005, w_039_136, w_052_061);
  or2  I058_007(w_058_007, w_021_031, w_026_098);
  not1 I058_010(w_058_010, w_021_108);
  or2  I058_012(w_058_012, w_027_001, w_022_035);
  nand2 I058_014(w_058_014, w_045_139, w_035_013);
  or2  I058_016(w_058_016, w_011_036, w_021_090);
  nand2 I058_017(w_058_017, w_042_131, w_019_004);
  not1 I058_020(w_058_020, w_018_037);
  not1 I058_021(w_058_021, w_033_027);
  nand2 I058_023(w_058_023, w_006_000, w_000_468);
  nand2 I058_024(w_058_024, w_014_228, w_052_039);
  or2  I058_025(w_058_025, w_044_062, w_001_003);
  or2  I058_027(w_058_027, w_033_011, w_051_101);
  and2 I058_031(w_058_031, w_022_109, w_005_179);
  and2 I058_032(w_058_032, w_013_037, w_033_037);
  or2  I058_034(w_058_034, w_055_002, w_002_020);
  nand2 I058_035(w_058_035, w_017_087, w_041_217);
  or2  I058_037(w_058_037, w_035_051, w_034_194);
  and2 I058_038(w_058_038, w_034_011, w_033_048);
  not1 I058_040(w_058_040, w_017_016);
  or2  I058_041(w_058_041, w_019_030, w_026_084);
  not1 I058_047(w_058_047, w_044_323);
  nand2 I058_048(w_058_048, w_004_408, w_047_350);
  nand2 I058_051(w_058_051, w_052_019, w_007_082);
  or2  I058_052(w_058_052, w_028_096, w_022_110);
  nand2 I058_056(w_058_056, w_022_095, w_035_018);
  and2 I058_058(w_058_058, w_019_048, w_014_215);
  not1 I058_059(w_058_059, w_049_139);
  and2 I058_062(w_058_062, w_033_012, w_047_050);
  nand2 I058_068(w_058_068, w_014_085, w_001_004);
  not1 I058_072(w_058_072, w_036_166);
  and2 I058_073(w_058_073, w_030_053, w_016_378);
  or2  I058_074(w_058_074, w_051_221, w_002_013);
  nand2 I058_075(w_058_075, w_004_193, w_010_153);
  not1 I058_076(w_058_076, w_023_016);
  and2 I058_079(w_058_079, w_004_232, w_022_033);
  nand2 I058_081(w_058_081, w_024_296, w_043_052);
  or2  I058_083(w_058_083, w_019_016, w_034_238);
  nand2 I058_084(w_058_084, w_001_002, w_057_060);
  not1 I058_086(w_058_086, w_054_057);
  nand2 I059_004(w_059_004, w_024_261, w_044_008);
  nand2 I059_018(w_059_018, w_046_174, w_002_018);
  or2  I059_025(w_059_025, w_058_086, w_027_257);
  not1 I059_028(w_059_028, w_008_150);
  or2  I059_032(w_059_032, w_057_006, w_007_270);
  or2  I059_041(w_059_041, w_054_013, w_003_004);
  nand2 I059_046(w_059_046, w_030_071, w_031_017);
  and2 I059_056(w_059_056, w_048_271, w_045_008);
  nand2 I059_063(w_059_063, w_027_295, w_006_000);
  or2  I059_072(w_059_072, w_027_004, w_019_000);
  nand2 I059_077(w_059_077, w_010_446, w_054_081);
  nand2 I059_095(w_059_095, w_013_066, w_024_072);
  or2  I059_100(w_059_100, w_000_165, w_031_043);
  and2 I059_120(w_059_120, w_006_000, w_057_008);
  not1 I059_121(w_059_121, w_033_030);
  and2 I059_133(w_059_133, w_052_027, w_014_034);
  nand2 I059_148(w_059_148, w_045_096, w_024_270);
  and2 I059_158(w_059_158, w_039_346, w_051_028);
  and2 I059_159(w_059_159, w_011_106, w_058_001);
  or2  I059_168(w_059_168, w_031_015, w_036_060);
  nand2 I059_169(w_059_169, w_032_008, w_000_310);
  not1 I059_191(w_059_191, w_033_028);
  and2 I059_195(w_059_195, w_004_166, w_013_220);
  or2  I059_199(w_059_199, w_006_000, w_036_113);
  not1 I059_211(w_059_211, w_034_088);
  and2 I059_216(w_059_216, w_013_177, w_033_055);
  and2 I059_217(w_059_217, w_044_074, w_033_002);
  not1 I059_223(w_059_223, w_033_003);
  not1 I059_233(w_059_233, w_002_013);
  or2  I059_237(w_059_237, w_022_161, w_006_000);
  not1 I059_255(w_059_255, w_047_134);
  and2 I059_256(w_059_256, w_044_021, w_034_037);
  and2 I059_260(w_059_260, w_029_113, w_025_359);
  nand2 I059_262(w_059_262, w_027_282, w_032_014);
  and2 I059_264(w_059_264, w_027_025, w_040_004);
  nand2 I059_267(w_059_267, w_052_009, w_031_004);
  nand2 I059_269(w_059_269, w_032_048, w_026_192);
  and2 I059_272(w_059_272, w_058_032, w_001_000);
  or2  I059_280(w_059_280, w_053_037, w_009_049);
  nand2 I059_284(w_059_284, w_057_003, w_049_185);
  or2  I059_288(w_059_288, w_037_010, w_042_193);
  and2 I059_293(w_059_293, w_039_108, w_053_027);
  nand2 I059_297(w_059_297, w_019_013, w_039_448);
  and2 I059_317(w_059_317, w_043_143, w_010_207);
  nand2 I059_318(w_059_318, w_047_293, w_035_040);
  nand2 I059_322(w_059_322, w_028_100, w_043_014);
  not1 I059_337(w_059_337, w_055_085);
  nand2 I059_341(w_059_341, w_056_048, w_043_198);
  not1 I059_344(w_059_344, w_048_085);
  not1 I059_346(w_059_346, w_055_005);
  not1 I059_348(w_059_348, w_026_175);
  or2  I059_351(w_059_351, w_027_075, w_024_189);
  and2 I059_358(w_059_358, w_014_011, w_034_084);
  nand2 I059_359(w_059_359, w_052_116, w_029_082);
  and2 I059_390(w_059_390, w_018_045, w_014_056);
  or2  I059_403(w_059_403, w_023_110, w_035_061);
  or2  I059_415(w_059_415, w_013_052, w_034_150);
  not1 I059_438(w_059_438, w_048_104);
  or2  I059_440(w_059_440, w_048_014, w_043_082);
  nand2 I059_444(w_059_444, w_032_073, w_058_074);
  or2  I059_445(w_059_445, w_006_000, w_041_024);
  nand2 I059_461(w_059_461, w_057_054, w_018_171);
  and2 I059_478(w_059_478, w_008_215, w_000_207);
  or2  I059_484(w_059_484, w_017_078, w_004_366);
  and2 I060_009(w_060_009, w_003_084, w_049_307);
  nand2 I060_010(w_060_010, w_015_117, w_003_020);
  or2  I060_011(w_060_011, w_018_084, w_054_014);
  not1 I060_017(w_060_017, w_048_055);
  nand2 I060_020(w_060_020, w_036_190, w_043_063);
  and2 I060_023(w_060_023, w_026_370, w_014_046);
  not1 I060_027(w_060_027, w_019_030);
  not1 I060_032(w_060_032, w_021_001);
  or2  I060_033(w_060_033, w_039_454, w_000_135);
  nand2 I060_040(w_060_040, w_041_222, w_011_337);
  nand2 I060_045(w_060_045, w_000_437, w_045_150);
  and2 I060_047(w_060_047, w_059_041, w_049_174);
  nand2 I060_049(w_060_049, w_057_057, w_040_004);
  or2  I060_050(w_060_050, w_056_010, w_022_076);
  nand2 I060_055(w_060_055, w_041_004, w_027_378);
  not1 I060_060(w_060_060, w_033_043);
  or2  I060_064(w_060_064, w_006_000, w_021_033);
  and2 I060_065(w_060_065, w_022_091, w_047_354);
  nand2 I060_089(w_060_089, w_032_041, w_035_041);
  not1 I060_096(w_060_096, w_048_216);
  and2 I060_111(w_060_111, w_055_065, w_038_086);
  not1 I060_117(w_060_117, w_049_201);
  and2 I060_124(w_060_124, w_054_205, w_006_000);
  not1 I060_125(w_060_125, w_002_001);
  or2  I060_135(w_060_135, w_008_067, w_042_270);
  or2  I060_142(w_060_142, w_031_055, w_022_127);
  and2 I060_144(w_060_144, w_021_005, w_008_320);
  or2  I060_153(w_060_153, w_053_022, w_005_184);
  or2  I060_166(w_060_166, w_047_329, w_021_029);
  and2 I060_174(w_060_174, w_007_043, w_036_044);
  and2 I060_179(w_060_179, w_042_126, w_057_035);
  and2 I060_184(w_060_184, w_050_192, w_037_049);
  or2  I060_187(w_060_187, w_047_318, w_019_026);
  and2 I060_194(w_060_194, w_020_136, w_013_190);
  not1 I060_220(w_060_220, w_036_095);
  and2 I060_226(w_060_226, w_019_025, w_026_073);
  not1 I060_242(w_060_242, w_020_091);
  not1 I060_260(w_060_260, w_035_017);
  and2 I060_267(w_060_267, w_023_269, w_057_034);
  nand2 I060_268(w_060_268, w_050_176, w_056_087);
  or2  I060_290(w_060_290, w_020_084, w_010_150);
  not1 I060_295(w_060_295, w_048_003);
  nand2 I060_303(w_060_303, w_052_086, w_046_145);
  not1 I060_315(w_060_315, w_013_146);
  not1 I060_322(w_060_322, w_023_000);
  not1 I060_334(w_060_334, w_046_218);
  nand2 I060_344(w_060_344, w_046_043, w_029_163);
  or2  I060_370(w_060_370, w_015_072, w_024_084);
  not1 I060_379(w_060_379, w_012_151);
  or2  I060_432(w_060_432, w_038_009, w_053_001);
  nand2 I061_000(w_061_000, w_009_027, w_030_140);
  or2  I061_008(w_061_008, w_024_036, w_058_052);
  or2  I061_014(w_061_014, w_052_006, w_048_054);
  and2 I061_023(w_061_023, w_011_178, w_040_000);
  not1 I061_024(w_061_024, w_022_051);
  or2  I061_025(w_061_025, w_017_000, w_025_423);
  nand2 I061_027(w_061_027, w_034_179, w_019_048);
  and2 I061_032(w_061_032, w_047_175, w_031_022);
  and2 I061_039(w_061_039, w_008_277, w_056_003);
  and2 I061_041(w_061_041, w_002_008, w_008_115);
  or2  I061_047(w_061_047, w_030_107, w_024_112);
  nand2 I061_050(w_061_050, w_036_169, w_018_141);
  or2  I061_062(w_061_062, w_046_107, w_018_134);
  or2  I061_066(w_061_066, w_053_013, w_049_174);
  or2  I061_072(w_061_072, w_042_058, w_052_008);
  and2 I061_094(w_061_094, w_031_003, w_006_000);
  not1 I061_114(w_061_114, w_019_018);
  nand2 I061_117(w_061_117, w_003_026, w_013_196);
  and2 I061_126(w_061_126, w_054_020, w_017_162);
  or2  I061_127(w_061_127, w_000_222, w_050_152);
  not1 I061_130(w_061_130, w_015_083);
  nand2 I061_144(w_061_144, w_038_041, w_022_065);
  nand2 I061_160(w_061_160, w_002_011, w_014_195);
  not1 I061_170(w_061_170, w_060_125);
  and2 I061_174(w_061_174, w_037_126, w_046_180);
  nand2 I061_178(w_061_178, w_002_021, w_009_122);
  or2  I061_190(w_061_190, w_033_048, w_030_098);
  not1 I061_199(w_061_199, w_027_228);
  nand2 I061_207(w_061_207, w_024_280, w_022_010);
  or2  I061_208(w_061_208, w_016_350, w_023_388);
  or2  I061_212(w_061_212, w_019_021, w_014_218);
  not1 I061_213(w_061_213, w_059_217);
  not1 I061_222(w_061_222, w_041_056);
  and2 I061_224(w_061_224, w_003_035, w_004_071);
  or2  I061_236(w_061_236, w_037_041, w_004_424);
  nand2 I061_242(w_061_242, w_010_163, w_049_297);
  nand2 I061_247(w_061_247, w_033_032, w_013_173);
  not1 I061_249(w_061_249, w_048_234);
  and2 I061_265(w_061_265, w_023_053, w_013_188);
  and2 I061_268(w_061_268, w_035_016, w_021_103);
  and2 I061_271(w_061_271, w_049_200, w_057_033);
  or2  I061_275(w_061_275, w_054_110, w_040_002);
  not1 I061_284(w_061_284, w_047_279);
  and2 I061_297(w_061_297, w_017_080, w_012_195);
  or2  I061_304(w_061_304, w_056_008, w_043_156);
  nand2 I061_309(w_061_309, w_013_129, w_009_225);
  not1 I061_314(w_061_314, w_007_372);
  nand2 I061_330(w_061_330, w_055_068, w_019_052);
  or2  I061_334(w_061_334, w_032_065, w_020_112);
  or2  I061_337(w_061_337, w_002_009, w_029_188);
  and2 I061_356(w_061_356, w_014_039, w_002_018);
  not1 I061_367(w_061_367, w_047_216);
  not1 I061_373(w_061_373, w_014_256);
  and2 I061_376(w_061_376, w_060_055, w_059_233);
  not1 I061_383(w_061_383, w_034_205);
  not1 I061_391(w_061_391, w_030_191);
  not1 I061_405(w_061_405, w_032_052);
  nand2 I061_406(w_061_406, w_017_055, w_007_266);
  not1 I061_412(w_061_412, w_032_122);
  and2 I061_421(w_061_421, w_004_271, w_031_001);
  not1 I062_000(w_062_000, w_059_032);
  nand2 I062_002(w_062_002, w_012_015, w_046_211);
  nand2 I062_003(w_062_003, w_011_166, w_061_297);
  and2 I062_004(w_062_004, w_053_002, w_040_003);
  and2 I062_005(w_062_005, w_041_255, w_038_086);
  nand2 I062_006(w_062_006, w_044_275, w_053_029);
  nand2 I062_007(w_062_007, w_051_164, w_060_174);
  not1 I062_008(w_062_008, w_055_049);
  or2  I062_009(w_062_009, w_037_117, w_034_075);
  nand2 I062_010(w_062_010, w_034_154, w_051_001);
  not1 I062_011(w_062_011, w_030_031);
  not1 I062_012(w_062_012, w_007_286);
  or2  I062_013(w_062_013, w_053_015, w_011_083);
  not1 I062_015(w_062_015, w_016_007);
  or2  I062_016(w_062_016, w_024_241, w_022_069);
  and2 I062_018(w_062_018, w_032_011, w_008_058);
  not1 I062_019(w_062_019, w_015_054);
  nand2 I062_020(w_062_020, w_004_020, w_034_281);
  not1 I063_003(w_063_003, w_013_116);
  not1 I063_005(w_063_005, w_023_334);
  and2 I063_006(w_063_006, w_051_018, w_059_148);
  and2 I063_010(w_063_010, w_057_012, w_004_277);
  or2  I063_011(w_063_011, w_037_032, w_061_000);
  not1 I063_013(w_063_013, w_008_130);
  or2  I063_020(w_063_020, w_033_010, w_061_405);
  nand2 I063_022(w_063_022, w_002_013, w_029_024);
  nand2 I063_024(w_063_024, w_058_073, w_000_310);
  nand2 I063_025(w_063_025, w_033_026, w_050_035);
  not1 I063_026(w_063_026, w_000_368);
  or2  I063_028(w_063_028, w_042_013, w_029_124);
  nand2 I063_030(w_063_030, w_013_227, w_035_024);
  nand2 I063_036(w_063_036, w_055_012, w_060_153);
  and2 I063_043(w_063_043, w_005_108, w_005_178);
  or2  I063_047(w_063_047, w_000_186, w_004_396);
  and2 I063_056(w_063_056, w_037_144, w_062_020);
  or2  I063_057(w_063_057, w_016_141, w_016_292);
  not1 I063_062(w_063_062, w_011_021);
  or2  I063_074(w_063_074, w_062_016, w_018_010);
  not1 I063_076(w_063_076, w_049_179);
  or2  I063_078(w_063_078, w_042_196, w_000_167);
  not1 I063_079(w_063_079, w_050_045);
  or2  I063_089(w_063_089, w_022_038, w_053_026);
  and2 I063_091(w_063_091, w_057_044, w_061_412);
  and2 I063_097(w_063_097, w_003_055, w_000_040);
  and2 I063_106(w_063_106, w_050_124, w_006_000);
  or2  I063_111(w_063_111, w_046_062, w_041_099);
  and2 I063_113(w_063_113, w_007_049, w_012_001);
  not1 I063_114(w_063_114, w_019_024);
  or2  I063_117(w_063_117, w_019_031, w_038_008);
  nand2 I063_118(w_063_118, w_017_014, w_010_224);
  nand2 I063_122(w_063_122, w_022_053, w_050_034);
  and2 I063_123(w_063_123, w_058_068, w_012_006);
  nand2 I063_139(w_063_139, w_034_027, w_003_036);
  or2  I063_141(w_063_141, w_029_189, w_014_011);
  and2 I063_150(w_063_150, w_010_416, w_041_130);
  nand2 I063_159(w_063_159, w_032_068, w_054_020);
  or2  I063_165(w_063_165, w_025_311, w_033_031);
  not1 I063_171(w_063_171, w_026_305);
  or2  I063_174(w_063_174, w_008_333, w_012_326);
  nand2 I063_179(w_063_179, w_045_099, w_006_000);
  not1 I063_197(w_063_197, w_037_140);
  nand2 I063_200(w_063_200, w_003_062, w_034_257);
  nand2 I063_206(w_063_206, w_029_243, w_002_010);
  nand2 I063_208(w_063_208, w_032_139, w_037_023);
  nand2 I063_218(w_063_218, w_047_151, w_006_000);
  or2  I063_222(w_063_222, w_027_183, w_051_218);
  nand2 I063_223(w_063_223, w_032_013, w_036_196);
  and2 I063_226(w_063_226, w_059_199, w_053_025);
  not1 I063_228(w_063_228, w_002_019);
  not1 I063_232(w_063_232, w_004_309);
  or2  I063_256(w_063_256, w_015_078, w_047_276);
  nand2 I064_000(w_064_000, w_018_213, w_031_011);
  or2  I064_001(w_064_001, w_004_408, w_045_231);
  not1 I064_002(w_064_002, w_063_150);
  or2  I064_003(w_064_003, w_035_088, w_011_142);
  nand2 I064_006(w_064_006, w_021_008, w_019_014);
  or2  I064_007(w_064_007, w_050_055, w_014_233);
  not1 I064_009(w_064_009, w_034_192);
  nand2 I064_011(w_064_011, w_043_215, w_033_018);
  or2  I064_014(w_064_014, w_024_086, w_003_039);
  or2  I064_015(w_064_015, w_058_059, w_037_052);
  or2  I064_017(w_064_017, w_028_082, w_020_028);
  or2  I064_018(w_064_018, w_054_044, w_014_084);
  not1 I064_020(w_064_020, w_008_026);
  and2 I064_022(w_064_022, w_028_058, w_017_100);
  or2  I064_023(w_064_023, w_000_214, w_015_080);
  and2 I064_024(w_064_024, w_035_034, w_026_036);
  nand2 I064_030(w_064_030, w_031_052, w_063_111);
  nand2 I064_031(w_064_031, w_028_174, w_018_160);
  and2 I064_032(w_064_032, w_044_070, w_000_152);
  and2 I064_034(w_064_034, w_059_415, w_011_124);
  and2 I064_035(w_064_035, w_057_020, w_019_009);
  not1 I064_039(w_064_039, w_041_006);
  or2  I064_044(w_064_044, w_050_039, w_060_290);
  nand2 I064_045(w_064_045, w_008_012, w_028_239);
  not1 I064_046(w_064_046, w_005_097);
  and2 I064_047(w_064_047, w_022_070, w_051_081);
  nand2 I064_052(w_064_052, w_009_192, w_011_317);
  and2 I064_053(w_064_053, w_030_175, w_045_119);
  and2 I064_058(w_064_058, w_051_008, w_019_037);
  not1 I064_060(w_064_060, w_009_103);
  nand2 I064_070(w_064_070, w_023_189, w_026_219);
  not1 I065_007(w_065_007, w_003_095);
  and2 I065_009(w_065_009, w_011_292, w_028_006);
  not1 I065_010(w_065_010, w_023_400);
  and2 I065_014(w_065_014, w_012_369, w_011_041);
  not1 I065_019(w_065_019, w_021_039);
  not1 I065_021(w_065_021, w_047_015);
  and2 I065_024(w_065_024, w_025_010, w_011_315);
  not1 I065_027(w_065_027, w_054_048);
  not1 I065_029(w_065_029, w_032_066);
  and2 I065_032(w_065_032, w_016_007, w_030_029);
  not1 I065_035(w_065_035, w_041_122);
  or2  I065_036(w_065_036, w_025_212, w_055_074);
  or2  I065_039(w_065_039, w_039_376, w_041_151);
  not1 I065_041(w_065_041, w_050_106);
  and2 I065_042(w_065_042, w_064_009, w_045_152);
  and2 I065_050(w_065_050, w_027_241, w_037_143);
  and2 I065_055(w_065_055, w_028_048, w_039_176);
  not1 I065_057(w_065_057, w_027_211);
  not1 I065_070(w_065_070, w_031_003);
  or2  I065_072(w_065_072, w_054_030, w_029_057);
  and2 I065_079(w_065_079, w_021_047, w_039_223);
  not1 I065_084(w_065_084, w_043_192);
  nand2 I065_093(w_065_093, w_044_110, w_046_040);
  and2 I065_094(w_065_094, w_035_001, w_012_239);
  nand2 I065_104(w_065_104, w_019_014, w_029_198);
  not1 I065_105(w_065_105, w_008_241);
  nand2 I065_109(w_065_109, w_012_214, w_050_014);
  not1 I065_110(w_065_110, w_055_055);
  or2  I065_112(w_065_112, w_038_022, w_037_119);
  or2  I065_121(w_065_121, w_051_154, w_042_120);
  not1 I065_124(w_065_124, w_063_010);
  nand2 I065_126(w_065_126, w_048_196, w_037_097);
  nand2 I065_133(w_065_133, w_053_023, w_064_000);
  not1 I065_136(w_065_136, w_041_167);
  not1 I065_151(w_065_151, w_009_191);
  or2  I065_158(w_065_158, w_063_118, w_047_405);
  and2 I065_159(w_065_159, w_026_105, w_005_170);
  or2  I065_182(w_065_182, w_013_094, w_024_187);
  not1 I065_185(w_065_185, w_007_100);
  not1 I065_191(w_065_191, w_048_074);
  nand2 I065_202(w_065_202, w_051_031, w_061_127);
  and2 I065_210(w_065_210, w_056_139, w_039_063);
  nand2 I065_214(w_065_214, w_023_335, w_034_036);
  not1 I065_219(w_065_219, w_021_021);
  or2  I066_002(w_066_002, w_021_090, w_059_120);
  nand2 I066_003(w_066_003, w_045_018, w_032_059);
  or2  I066_006(w_066_006, w_029_017, w_031_023);
  nand2 I066_013(w_066_013, w_062_012, w_035_077);
  not1 I066_014(w_066_014, w_045_193);
  not1 I066_031(w_066_031, w_051_130);
  not1 I066_036(w_066_036, w_022_085);
  or2  I066_038(w_066_038, w_041_260, w_040_006);
  or2  I066_060(w_066_060, w_005_058, w_043_161);
  nand2 I066_067(w_066_067, w_016_177, w_031_057);
  and2 I066_072(w_066_072, w_059_095, w_014_083);
  nand2 I066_074(w_066_074, w_057_018, w_064_070);
  not1 I066_080(w_066_080, w_019_014);
  or2  I066_097(w_066_097, w_033_056, w_031_019);
  not1 I066_098(w_066_098, w_001_001);
  and2 I066_108(w_066_108, w_039_109, w_013_054);
  nand2 I066_111(w_066_111, w_034_081, w_024_130);
  and2 I066_113(w_066_113, w_042_250, w_021_018);
  nand2 I066_116(w_066_116, w_051_110, w_016_052);
  not1 I066_117(w_066_117, w_009_192);
  nand2 I066_126(w_066_126, w_062_019, w_025_130);
  not1 I066_128(w_066_128, w_053_006);
  not1 I066_131(w_066_131, w_034_155);
  not1 I066_135(w_066_135, w_030_072);
  or2  I066_145(w_066_145, w_056_164, w_038_070);
  and2 I066_150(w_066_150, w_020_045, w_056_058);
  not1 I066_154(w_066_154, w_045_065);
  not1 I066_160(w_066_160, w_054_146);
  or2  I066_163(w_066_163, w_028_258, w_050_117);
  and2 I066_168(w_066_168, w_058_047, w_059_256);
  and2 I066_169(w_066_169, w_046_006, w_005_096);
  not1 I067_000(w_067_000, w_021_051);
  or2  I067_001(w_067_001, w_062_020, w_004_393);
  nand2 I067_003(w_067_003, w_004_468, w_001_003);
  and2 I067_004(w_067_004, w_047_253, w_025_276);
  and2 I067_006(w_067_006, w_046_084, w_007_101);
  and2 I067_007(w_067_007, w_028_004, w_056_109);
  not1 I067_008(w_067_008, w_060_242);
  or2  I067_009(w_067_009, w_065_009, w_053_002);
  and2 I067_014(w_067_014, w_007_002, w_016_087);
  and2 I067_015(w_067_015, w_060_166, w_023_373);
  or2  I067_016(w_067_016, w_038_022, w_009_134);
  nand2 I067_017(w_067_017, w_044_055, w_032_087);
  nand2 I067_020(w_067_020, w_015_113, w_062_000);
  nand2 I067_022(w_067_022, w_029_241, w_006_000);
  nand2 I067_023(w_067_023, w_056_015, w_044_258);
  and2 I067_025(w_067_025, w_039_463, w_019_028);
  or2  I067_026(w_067_026, w_037_042, w_059_269);
  or2  I067_029(w_067_029, w_035_018, w_055_051);
  nand2 I067_030(w_067_030, w_026_213, w_008_132);
  nand2 I067_031(w_067_031, w_047_330, w_024_190);
  nand2 I067_032(w_067_032, w_063_006, w_029_202);
  nand2 I067_033(w_067_033, w_066_113, w_017_005);
  or2  I067_035(w_067_035, w_040_003, w_024_053);
  and2 I067_036(w_067_036, w_060_027, w_034_097);
  nand2 I067_039(w_067_039, w_046_015, w_062_007);
  or2  I067_040(w_067_040, w_064_000, w_018_143);
  nand2 I067_044(w_067_044, w_010_076, w_022_036);
  and2 I067_045(w_067_045, w_056_036, w_025_159);
  nand2 I067_050(w_067_050, w_024_183, w_029_039);
  and2 I067_051(w_067_051, w_017_091, w_056_050);
  nand2 I067_055(w_067_055, w_048_019, w_057_054);
  nand2 I067_056(w_067_056, w_016_245, w_008_135);
  not1 I067_059(w_067_059, w_042_054);
  nand2 I067_060(w_067_060, w_054_172, w_060_011);
  and2 I067_061(w_067_061, w_036_077, w_063_005);
  and2 I067_062(w_067_062, w_054_034, w_058_010);
  not1 I068_000(w_068_000, w_021_093);
  or2  I068_002(w_068_002, w_025_320, w_043_242);
  nand2 I068_003(w_068_003, w_025_091, w_013_040);
  nand2 I068_006(w_068_006, w_002_019, w_015_001);
  not1 I068_009(w_068_009, w_011_055);
  and2 I068_011(w_068_011, w_022_052, w_019_001);
  not1 I068_012(w_068_012, w_020_113);
  or2  I068_014(w_068_014, w_044_169, w_057_005);
  not1 I068_016(w_068_016, w_028_000);
  nand2 I068_020(w_068_020, w_013_097, w_030_129);
  nand2 I068_022(w_068_022, w_036_141, w_051_078);
  and2 I068_025(w_068_025, w_022_140, w_003_072);
  not1 I068_032(w_068_032, w_053_023);
  or2  I068_036(w_068_036, w_025_014, w_010_041);
  or2  I068_040(w_068_040, w_031_042, w_034_219);
  nand2 I068_042(w_068_042, w_060_089, w_017_186);
  not1 I068_046(w_068_046, w_011_207);
  not1 I068_048(w_068_048, w_019_013);
  nand2 I068_051(w_068_051, w_012_359, w_000_376);
  and2 I068_053(w_068_053, w_039_153, w_027_028);
  not1 I068_055(w_068_055, w_017_050);
  not1 I068_058(w_068_058, w_005_224);
  nand2 I068_066(w_068_066, w_022_116, w_028_370);
  and2 I068_070(w_068_070, w_012_326, w_017_003);
  or2  I068_076(w_068_076, w_011_073, w_067_014);
  or2  I068_080(w_068_080, w_029_071, w_021_071);
  nand2 I068_087(w_068_087, w_011_189, w_028_070);
  or2  I068_090(w_068_090, w_065_042, w_015_096);
  not1 I068_093(w_068_093, w_002_011);
  nand2 I068_097(w_068_097, w_067_062, w_041_160);
  and2 I068_099(w_068_099, w_042_189, w_033_001);
  not1 I068_100(w_068_100, w_008_064);
  not1 I068_103(w_068_103, w_012_077);
  or2  I068_119(w_068_119, w_047_141, w_044_075);
  not1 I068_129(w_068_129, w_011_101);
  nand2 I068_136(w_068_136, w_052_116, w_034_108);
  and2 I068_138(w_068_138, w_020_038, w_037_036);
  nand2 I068_139(w_068_139, w_035_085, w_007_292);
  and2 I068_146(w_068_146, w_064_002, w_035_025);
  nand2 I068_149(w_068_149, w_046_182, w_050_052);
  or2  I068_150(w_068_150, w_006_000, w_003_100);
  or2  I068_151(w_068_151, w_035_075, w_005_123);
  not1 I068_155(w_068_155, w_038_074);
  nand2 I068_156(w_068_156, w_029_141, w_060_187);
  nand2 I069_000(w_069_000, w_037_057, w_057_016);
  or2  I069_006(w_069_006, w_052_004, w_045_090);
  nand2 I069_008(w_069_008, w_032_023, w_055_040);
  nand2 I069_009(w_069_009, w_039_448, w_027_299);
  and2 I069_012(w_069_012, w_040_006, w_027_215);
  not1 I069_015(w_069_015, w_063_079);
  not1 I069_017(w_069_017, w_057_053);
  nand2 I069_023(w_069_023, w_006_000, w_051_041);
  or2  I069_026(w_069_026, w_004_454, w_010_038);
  or2  I069_028(w_069_028, w_027_165, w_003_022);
  not1 I069_031(w_069_031, w_025_197);
  and2 I069_037(w_069_037, w_050_070, w_004_016);
  or2  I069_040(w_069_040, w_018_206, w_028_187);
  and2 I069_054(w_069_054, w_000_377, w_054_012);
  nand2 I069_058(w_069_058, w_008_091, w_052_051);
  or2  I069_063(w_069_063, w_047_013, w_048_147);
  not1 I069_064(w_069_064, w_010_337);
  not1 I069_065(w_069_065, w_022_092);
  and2 I069_068(w_069_068, w_019_028, w_061_222);
  nand2 I069_069(w_069_069, w_001_000, w_041_065);
  nand2 I069_085(w_069_085, w_026_087, w_013_109);
  not1 I069_089(w_069_089, w_024_040);
  not1 I069_091(w_069_091, w_050_002);
  or2  I069_097(w_069_097, w_038_041, w_036_229);
  not1 I069_106(w_069_106, w_041_113);
  nand2 I069_108(w_069_108, w_015_091, w_063_150);
  or2  I069_109(w_069_109, w_035_016, w_068_022);
  and2 I069_112(w_069_112, w_030_068, w_007_049);
  and2 I069_125(w_069_125, w_007_378, w_049_003);
  nand2 I069_128(w_069_128, w_029_247, w_059_444);
  and2 I069_130(w_069_130, w_040_002, w_030_137);
  nand2 I069_132(w_069_132, w_010_207, w_023_215);
  nand2 I069_134(w_069_134, w_065_214, w_038_020);
  not1 I069_144(w_069_144, w_044_326);
  nand2 I069_147(w_069_147, w_034_166, w_048_022);
  nand2 I069_149(w_069_149, w_003_058, w_038_046);
  not1 I069_157(w_069_157, w_027_438);
  or2  I069_158(w_069_158, w_059_358, w_064_030);
  and2 I069_160(w_069_160, w_019_021, w_060_033);
  or2  I069_165(w_069_165, w_003_024, w_021_058);
  and2 I070_000(w_070_000, w_040_000, w_045_182);
  and2 I070_002(w_070_002, w_046_179, w_052_036);
  and2 I070_003(w_070_003, w_039_483, w_061_114);
  and2 I070_004(w_070_004, w_018_156, w_029_242);
  or2  I070_005(w_070_005, w_041_064, w_040_006);
  and2 I070_007(w_070_007, w_019_043, w_019_002);
  or2  I070_009(w_070_009, w_043_111, w_022_032);
  and2 I070_017(w_070_017, w_020_031, w_046_183);
  and2 I070_018(w_070_018, w_022_033, w_026_372);
  not1 I070_022(w_070_022, w_043_065);
  and2 I070_024(w_070_024, w_044_127, w_048_109);
  or2  I070_031(w_070_031, w_030_160, w_068_099);
  or2  I070_032(w_070_032, w_017_045, w_013_063);
  and2 I070_034(w_070_034, w_006_000, w_014_101);
  nand2 I070_040(w_070_040, w_054_166, w_028_118);
  and2 I070_041(w_070_041, w_034_210, w_050_073);
  nand2 I070_042(w_070_042, w_012_266, w_067_009);
  and2 I070_046(w_070_046, w_024_133, w_012_314);
  or2  I070_047(w_070_047, w_060_020, w_025_282);
  or2  I070_048(w_070_048, w_042_234, w_049_219);
  not1 I070_053(w_070_053, w_032_195);
  not1 I070_055(w_070_055, w_008_263);
  not1 I070_058(w_070_058, w_055_068);
  nand2 I070_059(w_070_059, w_064_030, w_027_439);
  not1 I070_061(w_070_061, w_022_018);
  not1 I070_065(w_070_065, w_023_359);
  not1 I070_067(w_070_067, w_023_046);
  nand2 I070_068(w_070_068, w_022_003, w_023_373);
  or2  I070_070(w_070_070, w_017_179, w_024_115);
  nand2 I070_072(w_070_072, w_016_052, w_018_098);
  not1 I070_074(w_070_074, w_026_014);
  or2  I070_076(w_070_076, w_020_075, w_013_201);
  nand2 I070_079(w_070_079, w_058_005, w_000_306);
  or2  I070_081(w_070_081, w_046_132, w_029_243);
  not1 I070_084(w_070_084, w_054_063);
  not1 I070_085(w_070_085, w_026_003);
  not1 I070_087(w_070_087, w_017_108);
  or2  I070_090(w_070_090, w_036_043, w_067_033);
  and2 I070_091(w_070_091, w_052_018, w_009_233);
  and2 I070_094(w_070_094, w_062_019, w_005_187);
  not1 I070_095(w_070_095, w_019_046);
  and2 I070_099(w_070_099, w_069_112, w_013_055);
  not1 I071_004(w_071_004, w_013_034);
  and2 I071_005(w_071_005, w_008_207, w_023_034);
  or2  I071_010(w_071_010, w_062_008, w_030_080);
  and2 I071_020(w_071_020, w_046_028, w_044_259);
  nand2 I071_036(w_071_036, w_024_187, w_024_186);
  and2 I071_046(w_071_046, w_044_112, w_020_014);
  or2  I071_055(w_071_055, w_052_103, w_045_180);
  and2 I071_088(w_071_088, w_042_106, w_054_055);
  and2 I071_089(w_071_089, w_026_210, w_020_184);
  not1 I071_094(w_071_094, w_063_043);
  nand2 I071_104(w_071_104, w_062_012, w_028_096);
  not1 I071_116(w_071_116, w_051_003);
  and2 I071_122(w_071_122, w_015_034, w_068_046);
  not1 I071_147(w_071_147, w_019_038);
  or2  I071_148(w_071_148, w_006_000, w_070_003);
  or2  I071_156(w_071_156, w_055_031, w_017_003);
  not1 I071_158(w_071_158, w_049_030);
  nand2 I071_169(w_071_169, w_031_001, w_067_015);
  not1 I071_185(w_071_185, w_006_000);
  and2 I071_191(w_071_191, w_027_155, w_002_027);
  or2  I071_193(w_071_193, w_032_141, w_054_204);
  nand2 I071_205(w_071_205, w_046_008, w_056_020);
  nand2 I071_211(w_071_211, w_060_050, w_046_174);
  or2  I071_212(w_071_212, w_021_034, w_061_212);
  not1 I071_214(w_071_214, w_050_017);
  nand2 I071_225(w_071_225, w_046_122, w_044_210);
  or2  I071_235(w_071_235, w_063_030, w_065_191);
  or2  I071_270(w_071_270, w_056_149, w_048_103);
  nand2 I071_289(w_071_289, w_021_071, w_056_122);
  nand2 I071_294(w_071_294, w_022_010, w_032_172);
  nand2 I071_295(w_071_295, w_025_234, w_047_023);
  or2  I071_299(w_071_299, w_034_084, w_031_066);
  nand2 I071_311(w_071_311, w_041_059, w_015_013);
  or2  I071_321(w_071_321, w_026_049, w_035_027);
  and2 I071_347(w_071_347, w_064_070, w_003_039);
  and2 I071_348(w_071_348, w_046_185, w_029_149);
  and2 I071_352(w_071_352, w_044_281, w_030_016);
  or2  I071_354(w_071_354, w_050_175, w_038_032);
  nand2 I071_358(w_071_358, w_034_172, w_036_099);
  nand2 I071_362(w_071_362, w_057_024, w_055_022);
  and2 I071_367(w_071_367, w_030_055, w_011_082);
  or2  I071_389(w_071_389, w_054_070, w_037_081);
  or2  I071_394(w_071_394, w_059_025, w_051_003);
  not1 I071_395(w_071_395, w_063_089);
  or2  I071_410(w_071_410, w_057_015, w_058_068);
  and2 I072_006(w_072_006, w_070_099, w_039_354);
  or2  I072_007(w_072_007, w_024_140, w_028_047);
  and2 I072_008(w_072_008, w_020_059, w_071_348);
  or2  I072_011(w_072_011, w_018_215, w_005_000);
  nand2 I072_014(w_072_014, w_036_105, w_071_395);
  and2 I072_018(w_072_018, w_021_012, w_017_113);
  and2 I072_020(w_072_020, w_037_093, w_001_004);
  and2 I072_022(w_072_022, w_018_312, w_032_074);
  or2  I072_031(w_072_031, w_025_248, w_006_000);
  and2 I072_034(w_072_034, w_036_030, w_062_006);
  or2  I072_042(w_072_042, w_026_362, w_058_000);
  and2 I072_045(w_072_045, w_046_221, w_038_088);
  nand2 I072_048(w_072_048, w_050_003, w_012_284);
  and2 I072_050(w_072_050, w_021_099, w_000_260);
  nand2 I072_053(w_072_053, w_036_081, w_000_474);
  or2  I072_054(w_072_054, w_019_023, w_040_000);
  nand2 I072_058(w_072_058, w_067_007, w_017_080);
  not1 I072_064(w_072_064, w_027_120);
  not1 I072_065(w_072_065, w_044_245);
  or2  I072_067(w_072_067, w_064_047, w_009_036);
  not1 I072_068(w_072_068, w_016_082);
  or2  I072_073(w_072_073, w_004_386, w_025_318);
  and2 I072_074(w_072_074, w_043_103, w_005_125);
  and2 I072_075(w_072_075, w_017_061, w_004_059);
  nand2 I072_080(w_072_080, w_017_173, w_047_044);
  or2  I072_084(w_072_084, w_041_022, w_057_050);
  nand2 I072_086(w_072_086, w_023_051, w_050_112);
  and2 I072_088(w_072_088, w_046_178, w_068_032);
  not1 I072_096(w_072_096, w_038_058);
  or2  I072_097(w_072_097, w_053_016, w_025_026);
  and2 I072_100(w_072_100, w_031_016, w_069_000);
  or2  I072_102(w_072_102, w_005_073, w_008_139);
  not1 I072_104(w_072_104, w_003_018);
  not1 I073_001(w_073_001, w_069_089);
  not1 I073_007(w_073_007, w_044_184);
  not1 I073_009(w_073_009, w_032_074);
  nand2 I073_010(w_073_010, w_049_301, w_037_116);
  and2 I073_012(w_073_012, w_069_058, w_052_054);
  nand2 I073_014(w_073_014, w_012_363, w_033_051);
  not1 I073_016(w_073_016, w_045_094);
  nand2 I073_017(w_073_017, w_009_065, w_034_003);
  or2  I073_021(w_073_021, w_060_135, w_003_025);
  or2  I073_023(w_073_023, w_025_143, w_064_007);
  or2  I073_026(w_073_026, w_062_018, w_022_095);
  and2 I073_027(w_073_027, w_009_126, w_062_008);
  nand2 I073_028(w_073_028, w_008_179, w_025_220);
  and2 I073_036(w_073_036, w_061_271, w_019_018);
  nand2 I073_039(w_073_039, w_007_322, w_002_025);
  and2 I073_040(w_073_040, w_056_162, w_024_074);
  and2 I073_041(w_073_041, w_043_006, w_009_065);
  not1 I073_043(w_073_043, w_041_039);
  or2  I073_044(w_073_044, w_043_029, w_006_000);
  or2  I073_046(w_073_046, w_061_356, w_024_209);
  nand2 I073_069(w_073_069, w_015_054, w_014_028);
  or2  I073_072(w_073_072, w_008_120, w_033_019);
  or2  I073_074(w_073_074, w_056_046, w_004_433);
  or2  I073_078(w_073_078, w_041_154, w_030_066);
  and2 I073_099(w_073_099, w_007_381, w_003_004);
  or2  I073_101(w_073_101, w_029_031, w_000_267);
  and2 I073_111(w_073_111, w_011_177, w_053_026);
  and2 I073_117(w_073_117, w_022_049, w_019_016);
  or2  I073_123(w_073_123, w_057_052, w_066_128);
  and2 I073_125(w_073_125, w_071_046, w_000_281);
  nand2 I073_129(w_073_129, w_044_277, w_057_019);
  not1 I073_132(w_073_132, w_021_021);
  or2  I073_133(w_073_133, w_061_421, w_043_077);
  and2 I073_138(w_073_138, w_048_064, w_043_179);
  and2 I073_149(w_073_149, w_058_062, w_063_159);
  and2 I073_172(w_073_172, w_018_164, w_058_079);
  or2  I073_173(w_073_173, w_033_027, w_041_211);
  or2  I073_176(w_073_176, w_014_103, w_068_103);
  not1 I073_181(w_073_181, w_020_180);
  nand2 I073_187(w_073_187, w_043_233, w_038_070);
  and2 I073_189(w_073_189, w_040_000, w_046_010);
  not1 I073_191(w_073_191, w_029_189);
  or2  I073_218(w_073_218, w_067_050, w_049_137);
  or2  I073_222(w_073_222, w_018_118, w_041_114);
  nand2 I074_000(w_074_000, w_054_043, w_057_003);
  not1 I074_001(w_074_001, w_063_165);
  not1 I074_002(w_074_002, w_033_014);
  or2  I074_003(w_074_003, w_064_001, w_024_110);
  or2  I074_004(w_074_004, w_019_032, w_070_058);
  and2 I074_005(w_074_005, w_051_097, w_033_037);
  and2 I075_018(w_075_018, w_000_033, w_009_041);
  nand2 I075_020(w_075_020, w_003_077, w_013_103);
  or2  I075_021(w_075_021, w_057_057, w_003_052);
  and2 I075_022(w_075_022, w_019_049, w_067_006);
  nand2 I075_024(w_075_024, w_001_002, w_007_308);
  not1 I075_025(w_075_025, w_008_342);
  or2  I075_038(w_075_038, w_072_088, w_074_004);
  nand2 I075_040(w_075_040, w_073_099, w_067_026);
  nand2 I075_041(w_075_041, w_010_423, w_032_070);
  not1 I075_042(w_075_042, w_045_184);
  or2  I075_047(w_075_047, w_072_084, w_054_000);
  nand2 I075_053(w_075_053, w_011_294, w_016_367);
  nand2 I075_054(w_075_054, w_069_130, w_011_067);
  nand2 I075_056(w_075_056, w_046_161, w_036_181);
  not1 I075_067(w_075_067, w_023_100);
  not1 I075_070(w_075_070, w_014_093);
  nand2 I075_074(w_075_074, w_051_306, w_055_056);
  nand2 I075_080(w_075_080, w_015_072, w_004_091);
  not1 I075_081(w_075_081, w_059_348);
  or2  I075_084(w_075_084, w_017_117, w_050_073);
  and2 I075_087(w_075_087, w_050_060, w_053_016);
  nand2 I075_089(w_075_089, w_036_168, w_070_076);
  and2 I075_091(w_075_091, w_015_009, w_049_066);
  and2 I075_093(w_075_093, w_014_018, w_062_018);
  or2  I075_094(w_075_094, w_031_057, w_046_166);
  and2 I075_095(w_075_095, w_017_052, w_046_165);
  nand2 I075_099(w_075_099, w_029_201, w_020_106);
  not1 I075_100(w_075_100, w_025_150);
  not1 I075_103(w_075_103, w_052_048);
  not1 I075_109(w_075_109, w_011_021);
  not1 I075_113(w_075_113, w_029_225);
  not1 I075_118(w_075_118, w_035_077);
  not1 I075_121(w_075_121, w_046_125);
  nand2 I075_122(w_075_122, w_058_027, w_000_328);
  not1 I075_124(w_075_124, w_049_038);
  and2 I075_130(w_075_130, w_018_108, w_009_062);
  or2  I076_000(w_076_000, w_009_091, w_018_283);
  and2 I076_008(w_076_008, w_059_272, w_072_080);
  nand2 I076_009(w_076_009, w_045_171, w_039_272);
  and2 I076_011(w_076_011, w_007_063, w_067_035);
  nand2 I076_013(w_076_013, w_061_373, w_035_045);
  nand2 I076_018(w_076_018, w_017_122, w_023_138);
  nand2 I076_020(w_076_020, w_049_076, w_056_106);
  and2 I076_021(w_076_021, w_058_034, w_002_000);
  nand2 I076_023(w_076_023, w_046_006, w_068_048);
  not1 I076_026(w_076_026, w_067_017);
  or2  I076_029(w_076_029, w_009_143, w_017_019);
  not1 I076_031(w_076_031, w_040_002);
  or2  I076_033(w_076_033, w_035_048, w_036_204);
  or2  I076_039(w_076_039, w_006_000, w_051_028);
  nand2 I076_042(w_076_042, w_003_063, w_039_024);
  and2 I076_045(w_076_045, w_000_142, w_020_170);
  not1 I076_056(w_076_056, w_018_102);
  not1 I076_058(w_076_058, w_027_008);
  or2  I076_060(w_076_060, w_064_045, w_002_012);
  nand2 I076_062(w_076_062, w_007_208, w_011_097);
  or2  I076_065(w_076_065, w_021_022, w_000_232);
  not1 I076_068(w_076_068, w_031_050);
  or2  I076_069(w_076_069, w_039_394, w_025_287);
  or2  I076_070(w_076_070, w_031_045, w_054_040);
  or2  I076_075(w_076_075, w_039_204, w_018_031);
  nand2 I076_077(w_076_077, w_022_126, w_055_071);
  not1 I076_078(w_076_078, w_044_014);
  not1 I076_085(w_076_085, w_066_117);
  not1 I076_086(w_076_086, w_023_159);
  and2 I076_093(w_076_093, w_046_178, w_072_011);
  not1 I076_094(w_076_094, w_019_003);
  or2  I076_095(w_076_095, w_025_277, w_036_179);
  not1 I076_097(w_076_097, w_029_184);
  or2  I076_102(w_076_102, w_042_217, w_026_002);
  nand2 I076_104(w_076_104, w_005_093, w_012_002);
  or2  I076_107(w_076_107, w_001_005, w_043_059);
  not1 I076_115(w_076_115, w_012_250);
  not1 I077_012(w_077_012, w_068_040);
  not1 I077_024(w_077_024, w_013_057);
  or2  I077_029(w_077_029, w_051_124, w_068_040);
  or2  I077_037(w_077_037, w_021_018, w_059_351);
  or2  I077_038(w_077_038, w_051_033, w_058_025);
  or2  I077_052(w_077_052, w_046_122, w_024_144);
  and2 I077_053(w_077_053, w_045_008, w_013_001);
  not1 I077_057(w_077_057, w_061_144);
  not1 I077_061(w_077_061, w_030_030);
  or2  I077_083(w_077_083, w_038_009, w_044_013);
  and2 I077_085(w_077_085, w_016_139, w_053_014);
  nand2 I077_086(w_077_086, w_022_122, w_006_000);
  nand2 I077_099(w_077_099, w_010_427, w_020_113);
  or2  I077_101(w_077_101, w_072_022, w_005_105);
  or2  I077_104(w_077_104, w_002_019, w_009_014);
  and2 I077_109(w_077_109, w_048_190, w_016_371);
  not1 I077_113(w_077_113, w_050_128);
  nand2 I077_117(w_077_117, w_069_068, w_073_123);
  and2 I077_120(w_077_120, w_052_039, w_020_062);
  or2  I077_123(w_077_123, w_014_148, w_053_003);
  nand2 I077_125(w_077_125, w_039_104, w_064_011);
  and2 I077_135(w_077_135, w_033_005, w_020_001);
  not1 I077_142(w_077_142, w_005_042);
  or2  I077_148(w_077_148, w_067_031, w_047_256);
  or2  I077_153(w_077_153, w_002_007, w_036_006);
  or2  I077_156(w_077_156, w_033_054, w_032_004);
  nand2 I077_157(w_077_157, w_011_030, w_059_297);
  nand2 I077_162(w_077_162, w_071_367, w_008_054);
  and2 I077_164(w_077_164, w_037_149, w_014_196);
  or2  I077_174(w_077_174, w_072_104, w_020_150);
  not1 I077_184(w_077_184, w_016_189);
  not1 I077_185(w_077_185, w_051_151);
  or2  I077_191(w_077_191, w_075_070, w_062_012);
  not1 I077_201(w_077_201, w_054_064);
  and2 I077_236(w_077_236, w_023_277, w_045_118);
  not1 I077_246(w_077_246, w_046_148);
  or2  I078_000(w_078_000, w_063_179, w_054_100);
  and2 I078_001(w_078_001, w_030_128, w_067_029);
  or2  I078_002(w_078_002, w_065_057, w_055_005);
  not1 I078_006(w_078_006, w_003_005);
  not1 I078_011(w_078_011, w_034_152);
  not1 I078_012(w_078_012, w_003_076);
  nand2 I078_013(w_078_013, w_022_159, w_072_018);
  or2  I078_019(w_078_019, w_069_065, w_046_023);
  nand2 I078_028(w_078_028, w_070_079, w_061_062);
  not1 I078_032(w_078_032, w_063_171);
  or2  I078_041(w_078_041, w_038_012, w_050_007);
  or2  I078_050(w_078_050, w_034_084, w_052_084);
  or2  I078_053(w_078_053, w_040_005, w_069_125);
  not1 I078_055(w_078_055, w_067_031);
  nand2 I078_057(w_078_057, w_007_042, w_009_235);
  or2  I078_062(w_078_062, w_030_030, w_000_272);
  not1 I078_063(w_078_063, w_055_043);
  not1 I078_066(w_078_066, w_044_120);
  nand2 I078_067(w_078_067, w_045_094, w_006_000);
  not1 I078_071(w_078_071, w_058_001);
  and2 I078_074(w_078_074, w_073_041, w_009_143);
  not1 I078_078(w_078_078, w_071_156);
  nand2 I078_081(w_078_081, w_042_099, w_026_363);
  or2  I078_086(w_078_086, w_028_364, w_057_028);
  or2  I078_090(w_078_090, w_014_219, w_006_000);
  not1 I078_091(w_078_091, w_037_057);
  or2  I078_094(w_078_094, w_060_032, w_071_088);
  nand2 I078_099(w_078_099, w_008_138, w_075_022);
  nand2 I078_104(w_078_104, w_034_101, w_057_035);
  nand2 I078_107(w_078_107, w_008_040, w_061_247);
  or2  I078_116(w_078_116, w_065_079, w_012_341);
  and2 I078_117(w_078_117, w_024_222, w_023_235);
  and2 I078_123(w_078_123, w_023_353, w_021_036);
  nand2 I078_126(w_078_126, w_027_249, w_017_167);
  nand2 I078_136(w_078_136, w_028_237, w_047_274);
  and2 I078_142(w_078_142, w_068_009, w_066_031);
  not1 I078_143(w_078_143, w_017_101);
  or2  I078_144(w_078_144, w_009_007, w_061_008);
  or2  I078_160(w_078_160, w_032_026, w_009_120);
  and2 I078_161(w_078_161, w_055_035, w_039_421);
  not1 I078_163(w_078_163, w_004_295);
  or2  I078_164(w_078_164, w_051_041, w_063_057);
  or2  I079_007(w_079_007, w_057_021, w_055_028);
  not1 I079_013(w_079_013, w_041_168);
  and2 I079_020(w_079_020, w_041_007, w_012_181);
  or2  I079_021(w_079_021, w_036_147, w_058_035);
  nand2 I079_028(w_079_028, w_018_263, w_017_124);
  and2 I079_040(w_079_040, w_021_091, w_036_169);
  not1 I079_047(w_079_047, w_052_020);
  nand2 I079_065(w_079_065, w_004_061, w_034_058);
  or2  I079_133(w_079_133, w_053_033, w_015_045);
  nand2 I079_141(w_079_141, w_039_240, w_008_084);
  and2 I079_158(w_079_158, w_073_036, w_071_347);
  nand2 I079_170(w_079_170, w_014_119, w_068_003);
  not1 I079_181(w_079_181, w_009_220);
  nand2 I079_193(w_079_193, w_035_097, w_063_062);
  not1 I079_197(w_079_197, w_032_167);
  or2  I079_199(w_079_199, w_058_038, w_021_075);
  nand2 I079_219(w_079_219, w_008_254, w_056_047);
  nand2 I079_224(w_079_224, w_062_019, w_055_000);
  nand2 I079_235(w_079_235, w_052_048, w_013_001);
  and2 I079_237(w_079_237, w_061_304, w_032_098);
  not1 I079_247(w_079_247, w_008_134);
  or2  I079_256(w_079_256, w_032_058, w_062_011);
  or2  I079_257(w_079_257, w_016_319, w_046_180);
  and2 I079_267(w_079_267, w_011_115, w_057_059);
  or2  I079_304(w_079_304, w_017_126, w_018_151);
  or2  I079_320(w_079_320, w_037_029, w_014_017);
  and2 I079_328(w_079_328, w_035_094, w_027_196);
  not1 I079_342(w_079_342, w_035_004);
  not1 I079_362(w_079_362, w_050_039);
  or2  I079_401(w_079_401, w_024_127, w_076_060);
  or2  I079_402(w_079_402, w_012_290, w_055_086);
  and2 I079_407(w_079_407, w_058_072, w_046_208);
  and2 I079_422(w_079_422, w_045_039, w_069_132);
  not1 I079_432(w_079_432, w_048_012);
  not1 I079_434(w_079_434, w_076_023);
  not1 I079_452(w_079_452, w_041_052);
  nand2 I079_453(w_079_453, w_035_100, w_059_169);
  or2  I080_000(w_080_000, w_064_032, w_071_311);
  and2 I080_001(w_080_001, w_015_108, w_052_012);
  and2 I080_003(w_080_003, w_006_000, w_042_084);
  nand2 I080_004(w_080_004, w_027_443, w_006_000);
  not1 I080_005(w_080_005, w_048_303);
  and2 I080_007(w_080_007, w_018_301, w_071_169);
  and2 I080_009(w_080_009, w_056_054, w_070_070);
  or2  I080_011(w_080_011, w_070_004, w_003_048);
  or2  I080_012(w_080_012, w_004_203, w_056_063);
  and2 I080_013(w_080_013, w_024_166, w_037_075);
  and2 I080_014(w_080_014, w_006_000, w_057_002);
  not1 I080_015(w_080_015, w_026_104);
  not1 I080_016(w_080_016, w_048_128);
  not1 I080_017(w_080_017, w_076_069);
  or2  I080_018(w_080_018, w_060_267, w_008_053);
  nand2 I080_019(w_080_019, w_016_024, w_067_061);
  and2 I080_020(w_080_020, w_056_148, w_060_144);
  or2  I080_021(w_080_021, w_028_132, w_064_022);
  and2 I080_023(w_080_023, w_048_050, w_016_256);
  or2  I080_024(w_080_024, w_044_112, w_010_104);
  not1 I080_025(w_080_025, w_018_003);
  nand2 I080_028(w_080_028, w_033_016, w_039_367);
  nand2 I080_031(w_080_031, w_007_219, w_054_054);
  or2  I080_032(w_080_032, w_024_127, w_038_005);
  and2 I080_035(w_080_035, w_018_001, w_023_413);
  not1 I081_001(w_081_001, w_023_232);
  nand2 I081_003(w_081_003, w_045_229, w_046_115);
  nand2 I081_004(w_081_004, w_010_391, w_058_012);
  or2  I081_008(w_081_008, w_055_052, w_000_153);
  or2  I081_010(w_081_010, w_032_108, w_012_048);
  and2 I081_011(w_081_011, w_022_012, w_012_041);
  or2  I081_012(w_081_012, w_056_092, w_002_021);
  or2  I081_017(w_081_017, w_073_016, w_047_292);
  and2 I081_018(w_081_018, w_075_084, w_054_097);
  nand2 I081_020(w_081_020, w_035_066, w_030_146);
  nand2 I081_025(w_081_025, w_065_110, w_029_010);
  not1 I081_026(w_081_026, w_020_091);
  not1 I081_027(w_081_027, w_071_225);
  or2  I081_029(w_081_029, w_042_001, w_017_163);
  and2 I081_030(w_081_030, w_024_275, w_053_027);
  and2 I081_034(w_081_034, w_047_400, w_025_248);
  not1 I081_035(w_081_035, w_049_107);
  or2  I081_037(w_081_037, w_031_022, w_069_023);
  not1 I081_038(w_081_038, w_055_011);
  nand2 I081_039(w_081_039, w_064_031, w_057_022);
  nand2 I081_044(w_081_044, w_059_288, w_019_052);
  and2 I081_053(w_081_053, w_000_110, w_028_015);
  not1 I081_058(w_081_058, w_001_006);
  or2  I081_061(w_081_061, w_052_104, w_051_253);
  or2  I081_064(w_081_064, w_040_002, w_018_165);
  not1 I081_069(w_081_069, w_062_002);
  or2  I081_073(w_081_073, w_023_020, w_019_016);
  not1 I081_074(w_081_074, w_068_053);
  nand2 I081_082(w_081_082, w_008_020, w_016_380);
  and2 I081_083(w_081_083, w_001_005, w_032_077);
  and2 I081_084(w_081_084, w_045_106, w_046_134);
  not1 I081_087(w_081_087, w_042_110);
  or2  I081_088(w_081_088, w_069_160, w_008_132);
  not1 I081_089(w_081_089, w_040_000);
  not1 I081_090(w_081_090, w_041_072);
  and2 I082_000(w_082_000, w_023_072, w_026_355);
  or2  I082_002(w_082_002, w_037_020, w_017_084);
  nand2 I082_005(w_082_005, w_042_183, w_060_017);
  not1 I082_007(w_082_007, w_043_241);
  and2 I082_015(w_082_015, w_038_009, w_052_036);
  nand2 I082_018(w_082_018, w_060_268, w_042_200);
  or2  I082_027(w_082_027, w_080_035, w_003_028);
  and2 I082_032(w_082_032, w_021_022, w_043_092);
  not1 I082_038(w_082_038, w_048_117);
  or2  I082_039(w_082_039, w_078_053, w_049_025);
  or2  I082_053(w_082_053, w_073_039, w_072_058);
  and2 I082_059(w_082_059, w_051_197, w_047_336);
  and2 I082_088(w_082_088, w_045_199, w_022_131);
  or2  I082_101(w_082_101, w_018_234, w_072_100);
  not1 I082_103(w_082_103, w_050_174);
  and2 I082_106(w_082_106, w_041_038, w_041_132);
  and2 I082_113(w_082_113, w_067_039, w_043_037);
  and2 I082_122(w_082_122, w_010_438, w_025_293);
  not1 I082_125(w_082_125, w_031_027);
  nand2 I082_126(w_082_126, w_065_007, w_051_286);
  or2  I082_134(w_082_134, w_016_140, w_081_082);
  not1 I082_141(w_082_141, w_030_002);
  not1 I082_144(w_082_144, w_002_023);
  nand2 I082_158(w_082_158, w_026_266, w_070_059);
  or2  I082_188(w_082_188, w_078_142, w_044_146);
  not1 I082_196(w_082_196, w_076_045);
  or2  I082_197(w_082_197, w_021_083, w_001_005);
  nand2 I082_212(w_082_212, w_069_037, w_009_101);
  not1 I082_221(w_082_221, w_033_011);
  or2  I082_234(w_082_234, w_076_056, w_008_012);
  and2 I082_242(w_082_242, w_015_059, w_079_199);
  and2 I082_270(w_082_270, w_016_016, w_033_023);
  not1 I082_275(w_082_275, w_028_040);
  and2 I082_316(w_082_316, w_049_108, w_028_205);
  or2  I082_338(w_082_338, w_058_084, w_025_056);
  nand2 I082_339(w_082_341, w_080_021, w_082_340);
  or2  I082_340(w_082_342, w_082_341, w_017_104);
  not1 I082_341(w_082_343, w_082_342);
  or2  I082_342(w_082_344, w_082_343, w_057_048);
  not1 I082_343(w_082_345, w_082_344);
  and2 I082_344(w_082_340, w_007_357, w_082_345);
  nand2 I083_000(w_083_000, w_017_172, w_075_091);
  or2  I083_002(w_083_002, w_029_181, w_068_070);
  nand2 I083_003(w_083_003, w_065_041, w_004_001);
  not1 I083_004(w_083_004, w_040_003);
  nand2 I083_011(w_083_011, w_052_038, w_054_097);
  or2  I083_012(w_083_012, w_012_063, w_025_017);
  not1 I083_013(w_083_013, w_025_275);
  not1 I083_022(w_083_022, w_001_003);
  not1 I083_023(w_083_023, w_004_161);
  not1 I083_025(w_083_025, w_075_053);
  not1 I083_031(w_083_031, w_073_078);
  or2  I083_035(w_083_035, w_037_076, w_018_126);
  and2 I083_046(w_083_046, w_048_100, w_001_006);
  not1 I083_056(w_083_056, w_063_256);
  not1 I083_061(w_083_061, w_018_067);
  not1 I083_079(w_083_079, w_058_021);
  nand2 I083_083(w_083_083, w_053_011, w_000_255);
  not1 I083_084(w_083_084, w_077_057);
  or2  I083_090(w_083_090, w_014_095, w_067_025);
  nand2 I083_098(w_083_098, w_079_047, w_004_175);
  or2  I083_103(w_083_103, w_052_066, w_010_116);
  and2 I083_105(w_083_105, w_028_197, w_071_294);
  or2  I083_107(w_083_107, w_064_052, w_078_013);
  nand2 I083_108(w_083_108, w_078_063, w_082_158);
  nand2 I083_111(w_083_111, w_065_029, w_061_126);
  and2 I083_119(w_083_119, w_062_002, w_045_082);
  not1 I083_123(w_083_123, w_006_000);
  not1 I083_125(w_083_125, w_000_264);
  and2 I083_159(w_083_159, w_035_068, w_078_161);
  and2 I083_160(w_083_160, w_029_043, w_061_367);
  not1 I083_171(w_083_171, w_079_362);
  or2  I083_177(w_083_177, w_012_042, w_023_270);
  or2  I083_179(w_083_179, w_041_140, w_055_018);
  nand2 I083_188(w_083_188, w_027_194, w_019_050);
  not1 I083_195(w_083_195, w_063_097);
  nand2 I083_205(w_083_205, w_065_035, w_004_164);
  and2 I083_208(w_083_208, w_081_012, w_070_087);
  and2 I083_212(w_083_212, w_004_179, w_061_275);
  or2  I084_000(w_084_000, w_008_059, w_062_011);
  not1 I084_005(w_084_005, w_046_045);
  not1 I084_006(w_084_006, w_036_031);
  not1 I084_010(w_084_010, w_067_020);
  or2  I084_012(w_084_012, w_006_000, w_009_236);
  nand2 I084_020(w_084_020, w_071_321, w_035_090);
  not1 I084_026(w_084_026, w_077_109);
  or2  I084_030(w_084_030, w_026_137, w_005_149);
  and2 I084_031(w_084_031, w_082_039, w_064_047);
  nand2 I084_037(w_084_037, w_041_147, w_028_284);
  nand2 I084_051(w_084_051, w_070_067, w_038_051);
  or2  I084_053(w_084_053, w_051_056, w_064_022);
  and2 I084_055(w_084_055, w_021_066, w_004_269);
  not1 I084_062(w_084_062, w_069_109);
  nand2 I084_076(w_084_076, w_005_176, w_048_171);
  not1 I084_085(w_084_085, w_033_037);
  or2  I084_086(w_084_086, w_059_028, w_064_058);
  or2  I084_103(w_084_103, w_055_077, w_024_131);
  nand2 I084_111(w_084_111, w_018_136, w_017_050);
  or2  I084_113(w_084_113, w_024_153, w_080_031);
  and2 I084_114(w_084_114, w_054_073, w_038_011);
  or2  I084_122(w_084_122, w_000_444, w_076_031);
  not1 I084_132(w_084_132, w_076_093);
  not1 I084_136(w_084_136, w_019_046);
  not1 I084_137(w_084_137, w_034_138);
  not1 I084_163(w_084_163, w_030_091);
  or2  I084_176(w_084_176, w_056_137, w_061_391);
  and2 I084_201(w_084_201, w_076_042, w_018_278);
  not1 I084_207(w_084_207, w_022_028);
  nand2 I084_214(w_084_214, w_009_116, w_013_182);
  or2  I084_237(w_084_237, w_026_242, w_056_143);
  not1 I084_261(w_084_261, w_071_289);
  and2 I084_268(w_084_268, w_077_157, w_039_048);
  or2  I084_270(w_084_270, w_062_009, w_058_058);
  not1 I084_286(w_084_286, w_016_216);
  nand2 I084_288(w_084_288, w_028_379, w_026_242);
  nand2 I084_321(w_084_321, w_024_122, w_035_032);
  and2 I084_327(w_084_327, w_048_033, w_036_087);
  nand2 I084_337(w_084_337, w_065_039, w_065_094);
  and2 I084_342(w_084_342, w_024_214, w_078_160);
  and2 I085_002(w_085_002, w_025_014, w_009_090);
  not1 I085_017(w_085_017, w_033_031);
  or2  I085_021(w_085_021, w_019_022, w_054_068);
  not1 I085_027(w_085_027, w_007_007);
  not1 I085_036(w_085_036, w_076_011);
  not1 I085_044(w_085_044, w_054_210);
  nand2 I085_055(w_085_055, w_069_015, w_059_317);
  and2 I085_057(w_085_057, w_028_013, w_032_042);
  not1 I085_060(w_085_060, w_037_087);
  nand2 I085_065(w_085_065, w_021_040, w_022_043);
  nand2 I085_066(w_085_066, w_070_018, w_024_174);
  and2 I085_079(w_085_079, w_055_077, w_030_151);
  and2 I085_098(w_085_098, w_057_048, w_001_005);
  and2 I085_108(w_085_108, w_012_178, w_074_000);
  or2  I085_113(w_085_113, w_045_170, w_080_003);
  not1 I085_119(w_085_119, w_084_031);
  not1 I085_124(w_085_124, w_051_223);
  not1 I085_127(w_085_127, w_020_026);
  and2 I085_138(w_085_138, w_039_278, w_031_006);
  nand2 I085_139(w_085_139, w_042_145, w_062_011);
  nand2 I085_144(w_085_144, w_057_030, w_002_016);
  or2  I085_158(w_085_158, w_067_045, w_083_107);
  not1 I085_159(w_085_159, w_054_089);
  not1 I085_177(w_085_177, w_063_232);
  or2  I085_182(w_085_182, w_046_126, w_057_006);
  and2 I085_197(w_085_197, w_053_014, w_025_413);
  and2 I085_206(w_085_206, w_030_088, w_043_225);
  or2  I085_223(w_085_223, w_073_014, w_073_072);
  not1 I085_236(w_085_236, w_028_268);
  nand2 I085_244(w_085_244, w_062_002, w_015_074);
  or2  I085_246(w_085_246, w_035_046, w_071_148);
  not1 I086_001(w_086_001, w_045_114);
  not1 I086_007(w_086_007, w_068_076);
  not1 I086_010(w_086_010, w_015_068);
  nand2 I086_024(w_086_024, w_083_212, w_031_019);
  and2 I086_026(w_086_026, w_013_175, w_007_324);
  or2  I086_038(w_086_038, w_058_041, w_000_002);
  and2 I086_042(w_086_042, w_014_099, w_010_096);
  nand2 I086_043(w_086_043, w_073_028, w_017_166);
  or2  I086_047(w_086_047, w_072_014, w_076_058);
  and2 I086_052(w_086_052, w_016_044, w_005_145);
  and2 I086_055(w_086_055, w_036_027, w_063_174);
  nand2 I086_068(w_086_068, w_039_212, w_062_018);
  or2  I086_070(w_086_070, w_049_343, w_084_342);
  and2 I086_073(w_086_073, w_019_042, w_078_126);
  or2  I086_084(w_086_084, w_081_004, w_001_000);
  and2 I086_092(w_086_092, w_076_115, w_052_112);
  and2 I086_095(w_086_095, w_068_006, w_067_023);
  not1 I086_100(w_086_100, w_085_144);
  nand2 I086_102(w_086_102, w_072_086, w_006_000);
  not1 I086_103(w_086_103, w_077_101);
  or2  I086_107(w_086_107, w_056_046, w_009_020);
  and2 I086_120(w_086_120, w_057_004, w_030_138);
  nand2 I086_123(w_086_123, w_042_199, w_032_153);
  nand2 I086_133(w_086_133, w_059_158, w_005_110);
  and2 I086_140(w_086_140, w_027_006, w_051_119);
  nand2 I086_148(w_086_148, w_032_179, w_031_038);
  or2  I086_149(w_086_149, w_049_166, w_037_121);
  not1 I086_157(w_086_157, w_083_195);
  not1 I086_158(w_086_158, w_043_139);
  or2  I086_160(w_086_160, w_081_003, w_057_060);
  nand2 I086_161(w_086_161, w_051_159, w_081_058);
  not1 I086_165(w_086_165, w_007_072);
  or2  I086_188(w_086_188, w_055_036, w_050_155);
  nand2 I086_192(w_086_192, w_050_010, w_083_108);
  and2 I086_195(w_086_195, w_017_104, w_040_001);
  not1 I087_004(w_087_004, w_081_064);
  or2  I087_019(w_087_019, w_080_017, w_047_416);
  nand2 I087_027(w_087_027, w_004_251, w_053_035);
  not1 I087_038(w_087_038, w_028_221);
  and2 I087_039(w_087_039, w_004_339, w_070_042);
  or2  I087_061(w_087_061, w_003_029, w_084_288);
  nand2 I087_062(w_087_062, w_073_023, w_016_311);
  or2  I087_067(w_087_067, w_026_193, w_061_249);
  nand2 I087_074(w_087_074, w_020_042, w_058_024);
  or2  I087_082(w_087_082, w_003_019, w_004_282);
  nand2 I087_083(w_087_083, w_055_046, w_048_000);
  nand2 I087_104(w_087_104, w_028_266, w_062_007);
  or2  I087_130(w_087_130, w_038_007, w_081_090);
  and2 I087_138(w_087_138, w_059_159, w_062_020);
  nand2 I087_142(w_087_142, w_019_024, w_084_005);
  or2  I087_147(w_087_147, w_050_087, w_030_072);
  or2  I087_148(w_087_148, w_022_027, w_005_012);
  not1 I087_149(w_087_149, w_003_065);
  nand2 I087_178(w_087_178, w_015_082, w_037_075);
  and2 I087_188(w_087_188, w_034_048, w_081_083);
  or2  I087_217(w_087_217, w_078_107, w_043_230);
  nand2 I087_218(w_087_218, w_017_070, w_056_050);
  not1 I087_240(w_087_240, w_019_031);
  not1 I087_279(w_087_279, w_016_357);
  nand2 I087_281(w_087_281, w_048_209, w_015_116);
  and2 I087_314(w_087_314, w_043_007, w_000_031);
  or2  I087_322(w_087_322, w_071_116, w_040_005);
  not1 I088_012(w_088_012, w_066_002);
  or2  I088_021(w_088_021, w_052_040, w_036_118);
  not1 I088_030(w_088_030, w_069_134);
  not1 I088_031(w_088_031, w_065_109);
  and2 I088_041(w_088_041, w_064_039, w_086_188);
  and2 I088_061(w_088_061, w_058_047, w_042_206);
  not1 I088_107(w_088_107, w_003_036);
  and2 I088_119(w_088_119, w_046_007, w_046_040);
  nand2 I088_123(w_088_123, w_080_005, w_086_103);
  or2  I088_132(w_088_132, w_070_040, w_068_097);
  and2 I088_136(w_088_136, w_004_385, w_087_062);
  not1 I088_163(w_088_163, w_050_175);
  not1 I088_199(w_088_199, w_030_065);
  not1 I088_245(w_088_245, w_013_095);
  not1 I088_252(w_088_252, w_006_000);
  and2 I088_270(w_088_270, w_007_013, w_028_277);
  and2 I088_278(w_088_278, w_046_150, w_080_028);
  not1 I088_315(w_088_315, w_014_054);
  and2 I088_335(w_088_335, w_014_186, w_067_006);
  nand2 I088_336(w_088_336, w_077_117, w_013_192);
  nand2 I088_392(w_088_392, w_048_211, w_041_186);
  and2 I088_397(w_088_397, w_080_032, w_069_165);
  not1 I088_409(w_088_409, w_084_137);
  not1 I088_410(w_088_410, w_046_119);
  not1 I088_421(w_088_421, w_077_037);
  nand2 I088_435(w_088_435, w_039_224, w_053_019);
  not1 I088_445(w_088_445, w_063_025);
  not1 I088_453(w_088_455, w_088_454);
  or2  I088_454(w_088_456, w_088_455, w_088_471);
  not1 I088_455(w_088_454, w_088_456);
  nand2 I088_456(w_088_461, w_010_214, w_088_460);
  and2 I088_457(w_088_462, w_067_055, w_088_461);
  and2 I088_458(w_088_463, w_054_208, w_088_462);
  nand2 I088_459(w_088_464, w_088_463, w_047_234);
  nand2 I088_460(w_088_465, w_006_000, w_088_464);
  or2  I088_461(w_088_466, w_088_465, w_019_024);
  or2  I088_462(w_088_467, w_088_466, w_058_074);
  or2  I088_463(w_088_468, w_088_467, w_038_082);
  nand2 I088_464(w_088_469, w_073_043, w_088_468);
  not1 I088_465(w_088_460, w_088_456);
  and2 I088_466(w_088_471, w_026_204, w_088_469);
  nand2 I089_001(w_089_001, w_015_100, w_012_004);
  not1 I089_007(w_089_007, w_085_246);
  not1 I089_026(w_089_026, w_062_004);
  nand2 I089_031(w_089_031, w_076_018, w_074_004);
  nand2 I089_032(w_089_032, w_082_106, w_060_334);
  or2  I089_035(w_089_035, w_029_014, w_027_042);
  and2 I089_046(w_089_046, w_042_101, w_046_118);
  and2 I089_074(w_089_074, w_063_218, w_059_267);
  nand2 I089_090(w_089_090, w_030_078, w_021_083);
  or2  I089_092(w_089_092, w_059_216, w_010_408);
  and2 I089_096(w_089_096, w_081_089, w_060_040);
  not1 I089_101(w_089_101, w_047_174);
  or2  I089_103(w_089_103, w_000_374, w_084_321);
  not1 I089_120(w_089_120, w_069_147);
  not1 I089_138(w_089_138, w_023_269);
  not1 I089_180(w_089_180, w_017_101);
  and2 I089_189(w_089_189, w_085_127, w_083_025);
  and2 I089_193(w_089_193, w_077_153, w_024_112);
  or2  I089_217(w_089_217, w_020_119, w_088_392);
  nand2 I089_221(w_089_221, w_007_368, w_002_005);
  and2 I089_243(w_089_243, w_053_026, w_088_278);
  not1 I089_264(w_089_264, w_005_242);
  or2  I089_273(w_089_273, w_053_016, w_084_006);
  not1 I089_288(w_089_288, w_072_011);
  not1 I089_305(w_089_305, w_058_010);
  and2 I089_307(w_089_307, w_038_055, w_082_316);
  and2 I089_380(w_089_380, w_073_187, w_050_030);
  nand2 I089_400(w_089_400, w_062_000, w_011_329);
  not1 I089_404(w_089_404, w_036_094);
  or2  I089_416(w_089_416, w_087_149, w_074_003);
  and2 I089_429(w_089_429, w_076_107, w_020_107);
  or2  I089_431(w_089_431, w_076_008, w_041_033);
  and2 I089_442(w_089_442, w_058_023, w_016_018);
  and2 I090_012(w_090_012, w_030_176, w_083_123);
  or2  I090_017(w_090_017, w_009_185, w_047_045);
  or2  I090_019(w_090_019, w_065_112, w_005_028);
  and2 I090_064(w_090_064, w_015_075, w_076_075);
  and2 I090_068(w_090_068, w_010_052, w_046_023);
  and2 I090_076(w_090_076, w_014_135, w_057_046);
  and2 I090_079(w_090_079, w_020_164, w_015_006);
  and2 I090_087(w_090_087, w_058_081, w_063_197);
  nand2 I090_089(w_090_089, w_041_214, w_032_085);
  or2  I090_101(w_090_101, w_000_349, w_015_062);
  and2 I090_111(w_090_111, w_000_267, w_021_083);
  nand2 I090_120(w_090_120, w_048_029, w_031_024);
  not1 I090_128(w_090_128, w_007_315);
  not1 I090_139(w_090_139, w_071_212);
  not1 I090_141(w_090_141, w_025_172);
  and2 I090_163(w_090_163, w_061_213, w_008_276);
  and2 I090_177(w_090_177, w_028_216, w_013_127);
  nand2 I090_186(w_090_186, w_059_168, w_079_342);
  not1 I090_190(w_090_190, w_054_015);
  and2 I090_194(w_090_194, w_085_119, w_031_006);
  nand2 I090_215(w_090_215, w_024_128, w_057_010);
  not1 I090_221(w_090_221, w_049_273);
  nand2 I090_228(w_090_228, w_074_003, w_050_187);
  nand2 I090_249(w_090_249, w_016_002, w_039_309);
  or2  I090_256(w_090_256, w_029_001, w_014_010);
  and2 I090_262(w_090_262, w_060_017, w_085_138);
  not1 I090_281(w_090_281, w_027_313);
  not1 I090_283(w_090_283, w_028_009);
  or2  I090_287(w_090_287, w_039_040, w_047_316);
  not1 I090_288(w_090_288, w_025_262);
  nand2 I090_290(w_090_290, w_081_061, w_001_000);
  nand2 I090_298(w_090_298, w_065_070, w_018_076);
  and2 I090_301(w_090_301, w_002_018, w_075_021);
  and2 I090_317(w_090_317, w_081_011, w_043_143);
  nand2 I090_319(w_090_319, w_057_046, w_033_030);
  and2 I090_326(w_090_326, w_053_005, w_013_041);
  and2 I091_003(w_091_003, w_077_061, w_051_117);
  or2  I091_040(w_091_040, w_022_038, w_078_090);
  or2  I091_045(w_091_045, w_026_145, w_057_041);
  and2 I091_052(w_091_052, w_018_158, w_067_022);
  or2  I091_054(w_091_054, w_050_121, w_007_195);
  or2  I091_070(w_091_070, w_076_102, w_062_012);
  not1 I091_076(w_091_076, w_021_105);
  nand2 I091_077(w_091_077, w_046_044, w_023_081);
  not1 I091_109(w_091_109, w_031_058);
  and2 I091_123(w_091_123, w_062_015, w_064_034);
  nand2 I091_124(w_091_124, w_050_038, w_049_090);
  nand2 I091_135(w_091_135, w_041_000, w_076_000);
  and2 I091_152(w_091_152, w_047_415, w_073_074);
  not1 I091_168(w_091_168, w_045_004);
  nand2 I091_174(w_091_174, w_089_217, w_058_072);
  not1 I091_189(w_091_189, w_031_065);
  not1 I091_225(w_091_225, w_051_076);
  or2  I091_235(w_091_235, w_006_000, w_070_094);
  or2  I091_243(w_091_243, w_080_012, w_088_107);
  and2 I091_253(w_091_253, w_080_028, w_086_133);
  nand2 I091_254(w_091_254, w_083_013, w_043_064);
  and2 I091_258(w_091_258, w_065_084, w_046_097);
  not1 I091_260(w_091_260, w_070_058);
  not1 I091_264(w_091_264, w_015_065);
  nand2 I091_289(w_091_289, w_041_223, w_045_015);
  and2 I091_326(w_091_326, w_087_322, w_011_092);
  not1 I091_342(w_091_342, w_002_027);
  and2 I091_354(w_091_354, w_090_017, w_037_090);
  and2 I091_371(w_091_371, w_039_221, w_080_018);
  nand2 I091_411(w_091_411, w_047_258, w_021_007);
  not1 I091_417(w_091_417, w_078_012);
  or2  I092_005(w_092_005, w_029_222, w_038_099);
  or2  I092_009(w_092_009, w_049_266, w_070_024);
  not1 I092_014(w_092_014, w_081_020);
  nand2 I092_016(w_092_016, w_055_047, w_050_121);
  or2  I092_017(w_092_017, w_006_000, w_084_237);
  and2 I092_023(w_092_023, w_026_209, w_014_132);
  not1 I092_026(w_092_026, w_029_082);
  and2 I092_032(w_092_032, w_073_132, w_025_321);
  nand2 I092_033(w_092_033, w_054_003, w_006_000);
  or2  I092_035(w_092_035, w_005_078, w_018_157);
  not1 I092_038(w_092_038, w_003_088);
  and2 I092_045(w_092_045, w_006_000, w_062_010);
  or2  I092_049(w_092_049, w_057_060, w_072_007);
  nand2 I092_064(w_092_064, w_018_103, w_012_344);
  or2  I092_065(w_092_065, w_037_004, w_042_138);
  nand2 I092_068(w_092_068, w_076_039, w_087_038);
  or2  I092_073(w_092_073, w_024_285, w_022_069);
  or2  I092_074(w_092_074, w_082_122, w_016_262);
  and2 I092_076(w_092_076, w_026_326, w_079_402);
  not1 I092_085(w_092_085, w_090_089);
  and2 I092_087(w_092_087, w_025_045, w_046_138);
  and2 I092_094(w_092_094, w_040_004, w_070_024);
  not1 I092_107(w_092_107, w_090_256);
  or2  I092_109(w_092_109, w_067_059, w_011_268);
  and2 I092_112(w_092_112, w_008_011, w_057_005);
  not1 I092_123(w_092_123, w_042_142);
  nand2 I092_129(w_092_129, w_046_127, w_074_001);
  and2 I092_156(w_092_156, w_084_051, w_039_250);
  or2  I092_166(w_092_166, w_078_104, w_010_098);
  not1 I092_171(w_092_171, w_073_021);
  or2  I092_176(w_092_176, w_040_006, w_035_090);
  and2 I093_000(w_093_000, w_034_052, w_003_049);
  nand2 I093_004(w_093_004, w_088_410, w_045_177);
  and2 I093_009(w_093_009, w_023_233, w_073_069);
  not1 I093_018(w_093_018, w_065_019);
  or2  I093_024(w_093_024, w_092_087, w_084_020);
  not1 I093_034(w_093_034, w_001_000);
  nand2 I093_039(w_093_039, w_009_051, w_054_015);
  or2  I093_053(w_093_053, w_016_035, w_016_258);
  or2  I093_064(w_093_064, w_064_020, w_063_026);
  not1 I093_072(w_093_072, w_078_091);
  nand2 I093_095(w_093_095, w_030_144, w_076_008);
  nand2 I093_101(w_093_101, w_053_015, w_029_215);
  nand2 I093_107(w_093_107, w_085_057, w_087_130);
  and2 I093_110(w_093_110, w_013_023, w_075_118);
  or2  I093_111(w_093_111, w_041_186, w_009_192);
  not1 I093_115(w_093_115, w_045_216);
  and2 I093_143(w_093_143, w_053_034, w_005_073);
  and2 I093_152(w_093_152, w_017_186, w_069_054);
  or2  I093_161(w_093_161, w_086_043, w_040_002);
  nand2 I093_186(w_093_186, w_058_083, w_055_072);
  and2 I093_208(w_093_208, w_005_123, w_039_402);
  and2 I093_209(w_093_209, w_046_045, w_038_008);
  not1 I093_216(w_093_216, w_015_022);
  nand2 I093_246(w_093_246, w_059_255, w_012_309);
  and2 I093_258(w_093_258, w_039_077, w_054_005);
  nand2 I093_264(w_093_264, w_077_053, w_001_004);
  nand2 I093_266(w_093_266, w_038_013, w_011_073);
  and2 I093_269(w_093_269, w_015_047, w_007_047);
  or2  I093_272(w_093_272, w_089_180, w_047_231);
  not1 I093_276(w_093_276, w_001_002);
  and2 I093_281(w_093_281, w_081_010, w_032_176);
  not1 I093_293(w_093_293, w_071_354);
  not1 I093_295(w_093_295, w_034_247);
  or2  I093_318(w_093_318, w_090_177, w_017_035);
  and2 I093_329(w_093_329, w_058_056, w_062_019);
  not1 I093_346(w_093_346, w_076_078);
  or2  I093_348(w_093_348, w_081_018, w_044_297);
  nand2 I093_351(w_093_351, w_040_002, w_027_331);
  not1 I093_364(w_093_364, w_021_029);
  not1 I093_365(w_093_365, w_063_123);
  nand2 I093_371(w_093_371, w_023_404, w_055_047);
  and2 I093_378(w_093_378, w_048_207, w_014_208);
  and2 I093_425(w_093_427, w_093_426, w_018_293);
  nand2 I093_426(w_093_428, w_093_427, w_076_104);
  or2  I093_427(w_093_429, w_093_447, w_093_428);
  and2 I093_428(w_093_430, w_093_429, w_081_053);
  nand2 I093_429(w_093_426, w_043_071, w_093_430);
  nand2 I093_430(w_093_435, w_093_434, w_076_095);
  not1 I093_431(w_093_436, w_093_435);
  nand2 I093_432(w_093_437, w_093_436, w_067_030);
  nand2 I093_433(w_093_438, w_093_437, w_009_059);
  and2 I093_434(w_093_439, w_055_029, w_093_438);
  or2  I093_435(w_093_440, w_071_321, w_093_439);
  and2 I093_436(w_093_441, w_093_440, w_050_136);
  not1 I093_437(w_093_442, w_093_441);
  and2 I093_438(w_093_443, w_030_132, w_093_442);
  or2  I093_439(w_093_444, w_012_191, w_093_443);
  not1 I093_440(w_093_445, w_093_444);
  not1 I093_441(w_093_434, w_093_429);
  and2 I093_442(w_093_447, w_009_081, w_093_445);
  or2  I094_003(w_094_003, w_021_018, w_041_058);
  or2  I094_010(w_094_010, w_010_392, w_088_245);
  and2 I094_014(w_094_014, w_091_003, w_080_001);
  and2 I094_023(w_094_023, w_039_146, w_004_400);
  or2  I094_028(w_094_028, w_012_195, w_003_014);
  not1 I094_033(w_094_033, w_070_041);
  not1 I094_045(w_094_045, w_093_258);
  or2  I094_049(w_094_049, w_074_005, w_070_007);
  or2  I094_062(w_094_062, w_090_141, w_063_141);
  or2  I094_081(w_094_081, w_015_001, w_068_087);
  not1 I094_147(w_094_147, w_087_104);
  not1 I094_155(w_094_155, w_039_083);
  and2 I094_166(w_094_166, w_049_008, w_026_114);
  nand2 I094_171(w_094_171, w_055_002, w_040_001);
  or2  I094_199(w_094_199, w_020_104, w_011_115);
  and2 I094_229(w_094_229, w_004_228, w_082_234);
  or2  I094_319(w_094_319, w_003_047, w_070_002);
  nand2 I094_320(w_094_320, w_006_000, w_064_001);
  nand2 I094_357(w_094_357, w_016_014, w_084_268);
  or2  I094_393(w_094_393, w_046_062, w_047_368);
  nand2 I094_416(w_094_416, w_044_227, w_056_142);
  not1 I095_000(w_095_000, w_005_152);
  or2  I095_001(w_095_001, w_066_168, w_066_036);
  not1 I095_002(w_095_002, w_063_114);
  or2  I095_010(w_095_010, w_019_035, w_058_074);
  and2 I095_014(w_095_014, w_001_002, w_033_044);
  and2 I095_016(w_095_016, w_006_000, w_072_034);
  nand2 I095_017(w_095_017, w_068_093, w_021_049);
  not1 I095_023(w_095_023, w_036_127);
  or2  I095_026(w_095_026, w_038_077, w_011_021);
  or2  I095_030(w_095_030, w_080_001, w_060_009);
  or2  I095_036(w_095_036, w_088_252, w_071_410);
  not1 I095_037(w_095_037, w_015_089);
  and2 I095_038(w_095_038, w_013_220, w_061_309);
  or2  I095_044(w_095_044, w_079_432, w_060_117);
  or2  I095_048(w_095_048, w_016_030, w_077_156);
  or2  I095_049(w_095_049, w_003_043, w_038_008);
  nand2 I095_051(w_095_051, w_086_070, w_063_078);
  nand2 I095_052(w_095_052, w_086_123, w_093_161);
  not1 I095_058(w_095_058, w_010_064);
  and2 I095_061(w_095_061, w_043_022, w_058_048);
  and2 I095_064(w_095_064, w_038_082, w_008_053);
  or2  I095_066(w_095_066, w_067_055, w_045_004);
  not1 I095_067(w_095_067, w_079_256);
  and2 I095_073(w_095_073, w_002_024, w_071_104);
  not1 I095_080(w_095_080, w_019_019);
  nand2 I095_084(w_095_084, w_082_212, w_094_166);
  nand2 I095_089(w_095_089, w_029_124, w_038_009);
  or2  I095_091(w_095_091, w_091_045, w_031_048);
  and2 I095_094(w_095_094, w_000_401, w_032_142);
  or2  I095_099(w_095_099, w_045_104, w_024_148);
  or2  I096_004(w_096_004, w_051_146, w_091_371);
  or2  I096_009(w_096_009, w_004_400, w_004_190);
  and2 I096_010(w_096_010, w_010_328, w_046_021);
  not1 I096_017(w_096_017, w_064_053);
  or2  I096_018(w_096_018, w_033_039, w_021_075);
  or2  I096_020(w_096_020, w_036_155, w_023_083);
  not1 I096_022(w_096_022, w_013_222);
  and2 I096_024(w_096_024, w_048_285, w_048_021);
  nand2 I096_026(w_096_026, w_032_081, w_026_256);
  not1 I096_027(w_096_027, w_091_076);
  not1 I096_030(w_096_030, w_046_108);
  nand2 I096_033(w_096_033, w_072_007, w_087_019);
  and2 I096_038(w_096_038, w_074_000, w_029_215);
  and2 I096_039(w_096_039, w_027_108, w_003_079);
  not1 I096_046(w_096_046, w_002_020);
  or2  I096_054(w_096_054, w_007_072, w_086_158);
  or2  I096_059(w_096_059, w_063_208, w_065_050);
  or2  I096_086(w_096_086, w_093_186, w_061_207);
  not1 I096_095(w_096_095, w_014_173);
  or2  I096_102(w_096_102, w_032_041, w_007_178);
  or2  I096_106(w_096_106, w_053_031, w_089_431);
  and2 I096_127(w_096_127, w_042_177, w_000_252);
  not1 I096_134(w_096_134, w_080_016);
  and2 I096_136(w_096_136, w_029_111, w_059_461);
  or2  I096_145(w_096_145, w_094_393, w_083_046);
  not1 I096_146(w_096_146, w_010_208);
  and2 I096_147(w_096_147, w_063_036, w_056_053);
  and2 I096_150(w_096_150, w_002_004, w_037_126);
  nand2 I096_151(w_096_151, w_040_001, w_020_025);
  not1 I096_154(w_096_154, w_060_135);
  not1 I096_155(w_096_155, w_046_114);
  or2  I096_165(w_096_165, w_094_049, w_050_138);
  and2 I096_174(w_096_174, w_059_063, w_031_005);
  and2 I096_176(w_096_176, w_054_023, w_073_046);
  and2 I096_184(w_096_184, w_033_054, w_025_476);
  or2  I096_197(w_096_197, w_031_063, w_062_002);
  or2  I096_207(w_096_207, w_024_003, w_053_009);
  and2 I096_215(w_096_215, w_021_025, w_023_013);
  and2 I096_235(w_096_235, w_057_023, w_040_005);
  or2  I096_248(w_096_248, w_064_014, w_009_076);
  or2  I096_283(w_096_283, w_053_002, w_079_141);
  and2 I096_296(w_096_296, w_021_040, w_023_030);
  or2  I096_303(w_096_303, w_075_042, w_083_035);
  and2 I096_330(w_096_330, w_000_045, w_053_022);
  and2 I097_008(w_097_008, w_037_042, w_088_041);
  not1 I097_025(w_097_025, w_069_063);
  and2 I097_027(w_097_027, w_033_028, w_090_326);
  and2 I097_036(w_097_036, w_025_137, w_091_135);
  or2  I097_064(w_097_064, w_076_068, w_070_081);
  not1 I097_067(w_097_067, w_096_027);
  nand2 I097_070(w_097_070, w_037_011, w_041_075);
  or2  I097_092(w_097_092, w_012_245, w_004_160);
  or2  I097_097(w_097_097, w_043_071, w_004_244);
  not1 I097_111(w_097_111, w_042_092);
  or2  I097_114(w_097_114, w_034_191, w_093_152);
  and2 I097_125(w_097_125, w_055_028, w_019_006);
  nand2 I097_133(w_097_133, w_011_161, w_029_243);
  nand2 I097_139(w_097_139, w_016_068, w_068_103);
  nand2 I097_146(w_097_146, w_018_270, w_052_005);
  or2  I097_148(w_097_148, w_019_007, w_061_212);
  and2 I097_163(w_097_163, w_006_000, w_005_048);
  nand2 I097_164(w_097_164, w_071_122, w_049_000);
  not1 I097_165(w_097_165, w_028_073);
  and2 I097_167(w_097_167, w_062_005, w_023_150);
  nand2 I097_182(w_097_182, w_023_369, w_079_181);
  or2  I097_188(w_097_188, w_096_174, w_063_074);
  not1 I097_193(w_097_193, w_067_003);
  not1 I097_205(w_097_205, w_055_069);
  not1 I097_215(w_097_215, w_041_138);
  and2 I098_004(w_098_004, w_090_215, w_010_412);
  nand2 I098_005(w_098_005, w_003_047, w_029_097);
  and2 I098_006(w_098_006, w_093_295, w_035_041);
  not1 I098_008(w_098_008, w_042_067);
  and2 I098_009(w_098_009, w_048_233, w_047_089);
  or2  I098_010(w_098_010, w_062_010, w_014_240);
  or2  I098_011(w_098_011, w_060_010, w_087_027);
  nand2 I098_013(w_098_013, w_095_044, w_092_112);
  nand2 I098_014(w_098_014, w_018_175, w_021_000);
  or2  I098_015(w_098_015, w_013_162, w_006_000);
  nand2 I098_016(w_098_016, w_084_026, w_024_049);
  not1 I098_017(w_098_017, w_004_300);
  not1 I098_018(w_098_018, w_047_162);
  and2 I098_020(w_098_020, w_081_034, w_002_019);
  and2 I098_022(w_098_022, w_086_007, w_000_137);
  or2  I098_023(w_098_023, w_084_163, w_048_184);
  not1 I099_006(w_099_006, w_008_230);
  or2  I099_013(w_099_013, w_047_288, w_004_260);
  and2 I099_015(w_099_015, w_066_060, w_060_432);
  or2  I099_020(w_099_020, w_095_084, w_041_300);
  nand2 I099_022(w_099_022, w_012_339, w_008_053);
  nand2 I099_026(w_099_026, w_062_005, w_016_021);
  nand2 I099_037(w_099_037, w_027_389, w_050_182);
  and2 I099_038(w_099_038, w_063_091, w_036_028);
  not1 I099_043(w_099_043, w_002_004);
  nand2 I099_052(w_099_052, w_077_012, w_097_111);
  nand2 I099_054(w_099_054, w_097_036, w_034_154);
  or2  I099_056(w_099_056, w_049_380, w_063_011);
  and2 I099_059(w_099_059, w_096_197, w_068_025);
  not1 I099_075(w_099_075, w_060_295);
  and2 I099_088(w_099_088, w_076_086, w_010_035);
  nand2 I099_110(w_099_110, w_079_267, w_012_090);
  or2  I099_111(w_099_111, w_096_106, w_006_000);
  not1 I099_120(w_099_120, w_043_093);
  not1 I099_123(w_099_123, w_018_139);
  nand2 I099_150(w_099_150, w_006_000, w_034_077);
  nand2 I099_159(w_099_159, w_070_079, w_005_024);
  or2  I099_164(w_099_164, w_090_283, w_080_005);
  nand2 I099_180(w_099_180, w_037_043, w_080_031);
  and2 I099_181(w_099_181, w_071_358, w_065_158);
  and2 I099_196(w_099_196, w_026_007, w_022_093);
  or2  I099_223(w_099_223, w_037_014, w_059_337);
  not1 I099_226(w_099_226, w_021_070);
  not1 I099_244(w_099_244, w_036_131);
  or2  I099_267(w_099_267, w_034_193, w_031_008);
  or2  I099_271(w_099_271, w_077_142, w_048_137);
  nand2 I099_277(w_099_277, w_029_229, w_025_115);
  nand2 I100_003(w_100_003, w_079_422, w_050_187);
  and2 I100_035(w_100_035, w_063_003, w_081_074);
  nand2 I100_041(w_100_041, w_032_011, w_055_086);
  not1 I100_046(w_100_046, w_059_262);
  nand2 I100_062(w_100_062, w_096_033, w_051_010);
  nand2 I100_127(w_100_127, w_031_041, w_066_160);
  not1 I100_149(w_100_149, w_032_069);
  nand2 I100_157(w_100_157, w_034_177, w_079_197);
  not1 I100_163(w_100_163, w_041_185);
  and2 I100_179(w_100_179, w_022_036, w_011_112);
  not1 I100_180(w_100_180, w_045_201);
  nand2 I100_193(w_100_193, w_000_122, w_055_078);
  and2 I100_194(w_100_194, w_048_022, w_012_018);
  nand2 I100_215(w_100_215, w_059_403, w_075_100);
  and2 I100_219(w_100_219, w_004_081, w_072_031);
  and2 I100_230(w_100_230, w_051_124, w_052_098);
  or2  I100_231(w_100_231, w_017_071, w_096_046);
  and2 I100_258(w_100_258, w_030_078, w_093_266);
  nand2 I100_273(w_100_273, w_083_111, w_098_022);
  and2 I100_298(w_100_298, w_097_092, w_009_169);
  or2  I100_301(w_100_301, w_093_018, w_055_016);
  not1 I100_312(w_100_312, w_010_127);
  nand2 I100_402(w_100_402, w_060_322, w_007_269);
  and2 I101_001(w_101_001, w_074_000, w_024_018);
  nand2 I101_002(w_101_002, w_050_193, w_028_270);
  not1 I101_010(w_101_010, w_036_205);
  and2 I101_015(w_101_015, w_017_021, w_060_184);
  nand2 I101_019(w_101_019, w_001_004, w_064_060);
  nand2 I101_023(w_101_023, w_010_087, w_044_282);
  or2  I101_024(w_101_024, w_031_045, w_058_016);
  and2 I101_030(w_101_030, w_015_068, w_041_087);
  and2 I101_034(w_101_034, w_045_139, w_018_084);
  and2 I101_039(w_101_039, w_077_148, w_096_147);
  not1 I101_043(w_101_043, w_005_242);
  or2  I101_048(w_101_048, w_002_024, w_095_089);
  or2  I101_052(w_101_052, w_063_106, w_043_174);
  and2 I101_054(w_101_054, w_053_019, w_027_324);
  or2  I101_065(w_101_065, w_080_020, w_032_045);
  or2  I101_074(w_101_074, w_096_215, w_067_016);
  and2 I101_078(w_101_078, w_009_187, w_072_050);
  nand2 I101_099(w_101_099, w_100_231, w_096_095);
  and2 I101_101(w_101_101, w_068_006, w_057_027);
  and2 I101_105(w_101_105, w_076_104, w_036_157);
  or2  I101_106(w_101_106, w_002_020, w_051_210);
  and2 I101_126(w_101_126, w_097_114, w_091_243);
  not1 I101_128(w_101_128, w_003_087);
  nand2 I101_145(w_101_145, w_086_140, w_050_187);
  and2 I101_158(w_101_158, w_059_344, w_029_028);
  not1 I101_163(w_101_163, w_081_017);
  and2 I101_175(w_101_175, w_039_198, w_013_034);
  nand2 I101_186(w_101_186, w_096_095, w_090_249);
  or2  I101_201(w_101_201, w_096_303, w_077_052);
  or2  I101_225(w_101_225, w_098_004, w_014_046);
  or2  I101_249(w_101_249, w_036_108, w_000_231);
  not1 I101_254(w_101_254, w_095_067);
  not1 I101_270(w_101_270, w_071_020);
  nand2 I101_301(w_101_301, w_001_002, w_000_098);
  and2 I101_305(w_101_305, w_092_129, w_067_004);
  not1 I101_329(w_101_329, w_071_005);
  or2  I102_003(w_102_003, w_036_234, w_009_162);
  or2  I102_013(w_102_013, w_030_077, w_059_195);
  not1 I102_028(w_102_028, w_090_101);
  or2  I102_030(w_102_030, w_001_000, w_071_185);
  not1 I102_031(w_102_031, w_003_077);
  or2  I102_036(w_102_036, w_060_303, w_055_035);
  not1 I102_039(w_102_039, w_005_153);
  nand2 I102_044(w_102_044, w_057_051, w_044_157);
  and2 I102_047(w_102_047, w_076_033, w_004_447);
  and2 I102_059(w_102_059, w_056_068, w_002_008);
  and2 I102_071(w_102_071, w_059_438, w_046_151);
  nand2 I102_076(w_102_076, w_073_099, w_020_025);
  or2  I102_077(w_102_077, w_078_019, w_019_038);
  not1 I102_078(w_102_078, w_041_071);
  nand2 I102_079(w_102_079, w_053_013, w_054_051);
  not1 I102_080(w_102_080, w_021_058);
  not1 I102_083(w_102_083, w_075_095);
  not1 I102_087(w_102_087, w_025_350);
  nand2 I102_094(w_102_094, w_054_031, w_101_010);
  or2  I102_097(w_102_097, w_052_115, w_047_032);
  or2  I102_111(w_102_111, w_062_015, w_027_278);
  and2 I102_127(w_102_127, w_026_128, w_001_003);
  nand2 I102_129(w_102_129, w_011_334, w_053_027);
  not1 I102_131(w_102_131, w_010_042);
  or2  I102_147(w_102_147, w_016_002, w_026_013);
  and2 I102_149(w_102_149, w_055_074, w_059_237);
  nand2 I102_155(w_102_155, w_075_093, w_095_066);
  or2  I103_000(w_103_000, w_038_000, w_096_155);
  nand2 I103_001(w_103_001, w_017_180, w_095_048);
  not1 I103_002(w_103_002, w_083_159);
  or2  I103_003(w_103_003, w_047_278, w_093_216);
  and2 I103_004(w_103_004, w_067_031, w_034_252);
  not1 I103_005(w_103_005, w_088_409);
  nand2 I103_006(w_103_006, w_091_174, w_018_146);
  nand2 I103_007(w_103_007, w_056_058, w_044_161);
  not1 I103_008(w_103_008, w_062_013);
  nand2 I103_009(w_103_009, w_022_101, w_077_099);
  not1 I103_011(w_103_011, w_089_264);
  and2 I103_012(w_103_012, w_003_092, w_078_086);
  or2  I103_013(w_103_013, w_066_098, w_030_096);
  and2 I103_015(w_103_015, w_095_061, w_075_094);
  and2 I103_016(w_103_016, w_069_064, w_093_009);
  nand2 I103_017(w_103_017, w_095_036, w_021_104);
  not1 I103_018(w_103_018, w_011_026);
  or2  I104_002(w_104_002, w_050_184, w_011_011);
  and2 I104_007(w_104_007, w_044_074, w_048_001);
  and2 I104_014(w_104_014, w_039_080, w_033_021);
  or2  I104_022(w_104_022, w_062_011, w_036_227);
  or2  I104_026(w_104_026, w_082_242, w_073_138);
  not1 I104_031(w_104_031, w_002_016);
  nand2 I104_034(w_104_034, w_033_015, w_031_032);
  not1 I104_045(w_104_045, w_000_345);
  and2 I104_061(w_104_061, w_031_061, w_068_151);
  or2  I104_112(w_104_112, w_024_115, w_024_103);
  nand2 I104_129(w_104_129, w_099_037, w_030_150);
  not1 I104_192(w_104_192, w_026_036);
  or2  I104_223(w_104_223, w_091_253, w_055_033);
  or2  I104_260(w_104_260, w_034_195, w_035_046);
  and2 I104_263(w_104_263, w_089_103, w_078_001);
  or2  I104_301(w_104_301, w_030_080, w_081_037);
  nand2 I104_303(w_104_303, w_053_022, w_100_035);
  or2  I104_327(w_104_327, w_008_165, w_034_272);
  not1 I104_365(w_104_365, w_014_208);
  not1 I104_373(w_104_373, w_042_163);
  and2 I104_374(w_104_374, w_062_011, w_056_105);
  or2  I104_379(w_104_379, w_055_059, w_060_194);
  nand2 I104_385(w_104_385, w_024_150, w_100_230);
  nand2 I104_430(w_104_430, w_073_012, w_067_040);
  nand2 I105_001(w_105_001, w_099_043, w_017_116);
  and2 I105_012(w_105_012, w_091_342, w_049_002);
  and2 I105_026(w_105_026, w_049_173, w_056_118);
  or2  I105_033(w_105_033, w_002_011, w_023_376);
  and2 I105_035(w_105_035, w_009_133, w_095_001);
  or2  I105_041(w_105_041, w_002_022, w_036_143);
  or2  I105_047(w_105_047, w_048_284, w_046_170);
  and2 I105_051(w_105_051, w_072_086, w_098_009);
  or2  I105_057(w_105_057, w_087_130, w_024_074);
  not1 I105_077(w_105_077, w_079_007);
  nand2 I105_078(w_105_078, w_074_004, w_068_139);
  or2  I105_116(w_105_116, w_051_226, w_097_164);
  not1 I105_121(w_105_121, w_078_117);
  or2  I105_123(w_105_123, w_027_312, w_094_320);
  or2  I105_129(w_105_129, w_061_265, w_067_036);
  or2  I105_151(w_105_151, w_007_372, w_025_275);
  or2  I105_165(w_105_165, w_058_086, w_074_004);
  and2 I105_167(w_105_167, w_084_012, w_039_374);
  nand2 I105_177(w_105_177, w_015_043, w_055_045);
  and2 I105_192(w_105_192, w_054_083, w_087_218);
  or2  I105_231(w_105_231, w_029_184, w_005_110);
  and2 I105_246(w_105_246, w_010_134, w_012_065);
  or2  I105_248(w_105_248, w_088_021, w_007_063);
  not1 I105_293(w_105_293, w_080_016);
  or2  I105_297(w_105_297, w_047_154, w_057_054);
  and2 I105_317(w_105_317, w_008_218, w_033_003);
  and2 I105_382(w_105_382, w_073_009, w_026_230);
  not1 I105_426(w_105_426, w_027_337);
  or2  I106_003(w_106_003, w_049_323, w_071_214);
  and2 I106_007(w_106_007, w_015_112, w_079_020);
  and2 I106_010(w_106_010, w_067_020, w_043_218);
  nand2 I106_022(w_106_022, w_031_000, w_103_000);
  and2 I106_079(w_106_079, w_002_000, w_092_074);
  and2 I106_109(w_106_109, w_064_014, w_060_065);
  nand2 I106_146(w_106_146, w_086_026, w_086_157);
  and2 I106_164(w_106_164, w_058_031, w_050_204);
  and2 I106_168(w_106_168, w_097_188, w_011_257);
  not1 I106_176(w_106_176, w_057_037);
  and2 I106_184(w_106_184, w_043_217, w_062_012);
  nand2 I106_202(w_106_202, w_033_058, w_053_026);
  not1 I106_211(w_106_211, w_009_010);
  or2  I106_232(w_106_232, w_025_326, w_018_034);
  not1 I106_262(w_106_262, w_097_025);
  or2  I106_269(w_106_269, w_045_137, w_021_052);
  and2 I106_271(w_106_271, w_038_049, w_069_017);
  or2  I106_286(w_106_286, w_104_002, w_021_061);
  and2 I106_295(w_106_295, w_082_270, w_101_078);
  or2  I106_337(w_106_337, w_096_176, w_017_108);
  not1 I106_342(w_106_342, w_036_045);
  not1 I106_354(w_106_354, w_078_057);
  not1 I106_359(w_106_359, w_000_206);
  or2  I106_380(w_106_380, w_082_000, w_049_244);
  nand2 I106_395(w_106_395, w_095_002, w_030_091);
  nand2 I106_408(w_106_408, w_036_175, w_080_001);
  or2  I106_422(w_106_422, w_029_240, w_053_015);
  or2  I106_482(w_106_482, w_101_001, w_011_104);
  and2 I107_003(w_107_003, w_013_119, w_073_027);
  nand2 I107_010(w_107_010, w_035_037, w_021_027);
  or2  I107_013(w_107_013, w_106_109, w_006_000);
  not1 I107_021(w_107_021, w_019_053);
  and2 I107_022(w_107_022, w_104_045, w_047_174);
  not1 I107_023(w_107_023, w_004_105);
  nand2 I107_032(w_107_032, w_093_209, w_095_026);
  or2  I107_040(w_107_040, w_034_097, w_049_347);
  nand2 I107_041(w_107_041, w_091_054, w_074_003);
  or2  I107_043(w_107_043, w_004_019, w_065_032);
  or2  I107_045(w_107_045, w_007_322, w_056_048);
  not1 I107_046(w_107_046, w_094_171);
  or2  I107_047(w_107_047, w_075_018, w_032_103);
  not1 I107_056(w_107_056, w_058_076);
  or2  I107_057(w_107_057, w_005_106, w_023_172);
  and2 I107_058(w_107_058, w_052_033, w_073_101);
  and2 I107_061(w_107_061, w_102_031, w_105_231);
  or2  I107_067(w_107_067, w_048_118, w_019_006);
  or2  I107_068(w_107_068, w_018_144, w_079_028);
  nand2 I107_069(w_107_069, w_053_021, w_049_338);
  nand2 I108_000(w_108_000, w_016_011, w_006_000);
  nand2 I108_008(w_108_008, w_037_030, w_023_063);
  nand2 I108_010(w_108_010, w_031_056, w_013_132);
  not1 I108_011(w_108_011, w_083_083);
  not1 I108_017(w_108_017, w_009_011);
  and2 I108_019(w_108_019, w_083_061, w_041_291);
  or2  I108_023(w_108_023, w_030_066, w_031_020);
  or2  I108_024(w_108_024, w_099_164, w_050_102);
  or2  I108_025(w_108_025, w_035_006, w_066_080);
  not1 I108_028(w_108_028, w_063_057);
  nand2 I108_029(w_108_029, w_074_003, w_076_065);
  and2 I108_030(w_108_030, w_106_184, w_104_026);
  nand2 I108_032(w_108_032, w_055_076, w_093_095);
  or2  I108_036(w_108_036, w_056_074, w_053_015);
  and2 I108_038(w_108_038, w_069_157, w_100_046);
  nand2 I108_040(w_108_040, w_102_080, w_000_022);
  or2  I108_043(w_108_043, w_077_086, w_058_074);
  or2  I108_045(w_108_045, w_043_007, w_078_002);
  nand2 I108_046(w_108_046, w_001_005, w_050_047);
  and2 I108_050(w_108_050, w_083_205, w_020_107);
  nand2 I108_056(w_108_056, w_090_301, w_027_211);
  not1 I109_000(w_109_000, w_097_125);
  or2  I109_001(w_109_001, w_021_015, w_051_107);
  not1 I110_005(w_110_005, w_108_023);
  and2 I110_007(w_110_007, w_070_005, w_091_124);
  not1 I110_008(w_110_008, w_075_094);
  and2 I110_020(w_110_020, w_009_142, w_024_284);
  and2 I110_027(w_110_027, w_059_077, w_026_060);
  not1 I110_034(w_110_034, w_014_152);
  or2  I110_035(w_110_035, w_017_043, w_058_052);
  or2  I110_041(w_110_041, w_032_082, w_003_067);
  and2 I110_049(w_110_049, w_033_035, w_000_167);
  or2  I110_051(w_110_051, w_088_136, w_029_184);
  or2  I110_060(w_110_060, w_098_014, w_101_101);
  and2 I110_094(w_110_094, w_021_102, w_062_012);
  nand2 I110_095(w_110_095, w_037_065, w_057_039);
  or2  I110_132(w_110_132, w_078_099, w_056_054);
  nand2 I110_142(w_110_142, w_044_091, w_025_285);
  not1 I110_149(w_110_149, w_090_064);
  or2  I110_156(w_110_156, w_096_102, w_031_062);
  and2 I110_161(w_110_161, w_020_065, w_019_032);
  nand2 I110_172(w_110_172, w_041_139, w_044_171);
  or2  I110_193(w_110_193, w_093_348, w_089_429);
  and2 I110_194(w_110_194, w_048_304, w_022_058);
  or2  I110_210(w_110_210, w_022_000, w_076_070);
  nand2 I111_001(w_111_001, w_017_056, w_047_196);
  or2  I111_005(w_111_005, w_108_010, w_004_246);
  not1 I111_007(w_111_007, w_070_091);
  not1 I111_014(w_111_014, w_013_195);
  and2 I111_015(w_111_015, w_075_080, w_090_120);
  and2 I111_017(w_111_017, w_062_003, w_021_020);
  or2  I111_020(w_111_020, w_103_013, w_051_165);
  not1 I111_024(w_111_024, w_093_378);
  or2  I111_028(w_111_028, w_089_035, w_050_017);
  and2 I111_030(w_111_030, w_016_149, w_052_016);
  not1 I111_036(w_111_036, w_104_022);
  nand2 I111_037(w_111_037, w_045_038, w_032_158);
  and2 I111_047(w_111_047, w_015_061, w_033_003);
  nand2 I111_048(w_111_048, w_023_009, w_033_019);
  nand2 I111_055(w_111_055, w_099_120, w_009_132);
  not1 I111_061(w_111_061, w_092_085);
  or2  I111_066(w_111_066, w_088_132, w_069_015);
  or2  I111_069(w_111_069, w_031_048, w_065_112);
  not1 I111_081(w_111_081, w_027_404);
  or2  I111_087(w_111_087, w_026_004, w_019_020);
  or2  I111_088(w_111_088, w_083_160, w_016_028);
  and2 I112_017(w_112_017, w_037_130, w_023_075);
  or2  I112_020(w_112_020, w_012_238, w_071_158);
  nand2 I112_028(w_112_028, w_004_345, w_080_019);
  not1 I112_033(w_112_033, w_064_006);
  nand2 I112_035(w_112_035, w_110_005, w_083_022);
  nand2 I112_050(w_112_050, w_012_175, w_109_001);
  or2  I112_053(w_112_053, w_111_017, w_093_371);
  or2  I112_071(w_112_071, w_001_005, w_056_138);
  and2 I112_073(w_112_073, w_083_000, w_032_065);
  and2 I112_074(w_112_074, w_109_001, w_055_053);
  or2  I112_078(w_112_078, w_104_022, w_020_075);
  not1 I112_081(w_112_081, w_101_030);
  or2  I112_098(w_112_098, w_041_006, w_021_081);
  not1 I112_103(w_112_103, w_032_035);
  and2 I112_105(w_112_105, w_006_000, w_061_023);
  nand2 I112_108(w_112_108, w_109_001, w_077_038);
  and2 I112_131(w_112_131, w_020_012, w_052_101);
  or2  I112_142(w_112_142, w_036_261, w_008_296);
  nand2 I112_150(w_112_150, w_054_115, w_013_006);
  or2  I112_156(w_112_156, w_021_043, w_068_138);
  or2  I112_184(w_112_184, w_023_059, w_105_123);
  or2  I112_212(w_112_212, w_111_036, w_040_000);
  not1 I112_232(w_112_232, w_032_061);
  or2  I112_304(w_112_304, w_066_116, w_090_076);
  nand2 I112_363(w_112_363, w_075_130, w_033_010);
  or2  I113_002(w_113_002, w_007_382, w_101_015);
  or2  I113_007(w_113_007, w_002_018, w_032_106);
  nand2 I113_010(w_113_010, w_034_058, w_099_052);
  or2  I113_014(w_113_014, w_105_151, w_052_049);
  or2  I113_020(w_113_020, w_002_023, w_065_126);
  and2 I113_030(w_113_030, w_086_192, w_014_182);
  not1 I113_035(w_113_035, w_099_026);
  and2 I113_039(w_113_039, w_005_091, w_069_158);
  nand2 I113_041(w_113_041, w_080_007, w_066_013);
  nand2 I113_042(w_113_042, w_098_022, w_019_025);
  not1 I113_045(w_113_045, w_084_085);
  not1 I113_048(w_113_048, w_096_026);
  or2  I113_052(w_113_052, w_084_103, w_070_087);
  or2  I113_056(w_113_056, w_003_023, w_084_085);
  and2 I113_059(w_113_059, w_038_079, w_085_177);
  and2 I113_062(w_113_062, w_035_056, w_010_282);
  and2 I113_066(w_113_066, w_027_184, w_037_060);
  and2 I113_072(w_113_072, w_073_007, w_102_039);
  and2 I113_075(w_113_075, w_033_035, w_084_000);
  not1 I114_001(w_114_001, w_105_177);
  or2  I114_015(w_114_015, w_057_054, w_005_112);
  and2 I114_022(w_114_022, w_052_012, w_102_047);
  and2 I114_027(w_114_027, w_097_165, w_089_026);
  or2  I114_038(w_114_038, w_080_005, w_031_008);
  not1 I114_040(w_114_040, w_002_016);
  not1 I114_048(w_114_048, w_105_192);
  or2  I114_050(w_114_050, w_034_059, w_016_249);
  not1 I114_057(w_114_057, w_085_236);
  not1 I114_058(w_114_058, w_086_148);
  or2  I114_077(w_114_077, w_107_067, w_065_055);
  and2 I114_080(w_114_080, w_040_005, w_047_228);
  or2  I114_092(w_114_092, w_099_059, w_068_156);
  or2  I114_098(w_114_098, w_050_022, w_006_000);
  or2  I114_102(w_114_102, w_092_064, w_111_014);
  or2  I114_115(w_114_115, w_082_059, w_006_000);
  nand2 I114_146(w_114_146, w_071_094, w_010_051);
  nand2 I114_153(w_114_153, w_092_016, w_055_035);
  and2 I114_159(w_114_159, w_066_145, w_028_149);
  not1 I114_181(w_114_181, w_054_118);
  or2  I114_187(w_114_187, w_090_290, w_053_034);
  nand2 I114_188(w_114_188, w_050_138, w_088_336);
  and2 I114_192(w_114_192, w_028_009, w_005_212);
  not1 I114_195(w_114_195, w_095_023);
  nand2 I114_208(w_114_208, w_039_177, w_041_025);
  not1 I114_237(w_114_237, w_036_095);
  and2 I114_265(w_114_267, w_114_266, w_085_060);
  nand2 I114_266(w_114_268, w_114_267, w_113_062);
  not1 I114_267(w_114_269, w_114_268);
  and2 I114_268(w_114_270, w_114_269, w_055_001);
  and2 I114_269(w_114_271, w_027_444, w_114_270);
  and2 I114_270(w_114_272, w_110_132, w_114_271);
  not1 I114_271(w_114_273, w_114_272);
  or2  I114_272(w_114_274, w_096_038, w_114_273);
  nand2 I114_273(w_114_275, w_078_123, w_114_274);
  nand2 I114_274(w_114_276, w_114_289, w_114_275);
  nand2 I114_275(w_114_266, w_061_314, w_114_276);
  nand2 I114_276(w_114_281, w_114_280, w_068_080);
  or2  I114_277(w_114_282, w_060_379, w_114_281);
  and2 I114_278(w_114_283, w_035_079, w_114_282);
  not1 I114_279(w_114_284, w_114_283);
  or2  I114_280(w_114_285, w_050_146, w_114_284);
  or2  I114_281(w_114_286, w_114_285, w_073_189);
  or2  I114_282(w_114_287, w_012_020, w_114_286);
  not1 I114_283(w_114_280, w_114_276);
  and2 I114_284(w_114_289, w_074_005, w_114_287);
  or2  I115_031(w_115_031, w_009_158, w_011_041);
  not1 I115_032(w_115_032, w_084_201);
  not1 I115_037(w_115_037, w_047_286);
  or2  I115_095(w_115_095, w_046_032, w_025_029);
  and2 I115_131(w_115_131, w_008_132, w_003_075);
  not1 I115_164(w_115_164, w_073_010);
  and2 I115_171(w_115_171, w_105_051, w_042_067);
  and2 I115_174(w_115_174, w_027_268, w_088_123);
  or2  I115_185(w_115_185, w_023_284, w_006_000);
  not1 I115_195(w_115_195, w_070_048);
  nand2 I115_203(w_115_203, w_100_127, w_058_040);
  and2 I115_212(w_115_212, w_030_053, w_034_089);
  or2  I115_242(w_115_242, w_072_102, w_038_014);
  or2  I115_247(w_115_247, w_052_104, w_113_007);
  or2  I115_308(w_115_308, w_030_059, w_001_003);
  and2 I115_314(w_115_314, w_083_000, w_021_025);
  nand2 I115_320(w_115_320, w_027_341, w_044_108);
  or2  I115_330(w_115_330, w_093_034, w_032_051);
  and2 I115_346(w_115_346, w_053_009, w_005_064);
  or2  I115_379(w_115_379, w_077_117, w_010_344);
  and2 I115_423(w_115_423, w_028_201, w_099_196);
  nand2 I115_424(w_115_424, w_064_015, w_005_096);
  and2 I115_465(w_114_278, w_060_124, w_114_266);
  or2  I116_022(w_116_022, w_033_003, w_043_037);
  nand2 I116_023(w_116_023, w_108_000, w_082_005);
  nand2 I116_026(w_116_026, w_053_002, w_111_047);
  or2  I116_028(w_116_028, w_021_049, w_062_005);
  nand2 I116_029(w_116_029, w_097_067, w_010_353);
  nand2 I116_037(w_116_037, w_057_056, w_086_092);
  or2  I116_038(w_116_038, w_031_001, w_068_146);
  not1 I116_054(w_116_054, w_016_381);
  nand2 I116_059(w_116_059, w_025_325, w_009_045);
  or2  I116_094(w_116_094, w_054_042, w_077_191);
  or2  I116_100(w_116_100, w_089_221, w_083_046);
  and2 I116_108(w_116_108, w_058_079, w_081_044);
  and2 I116_116(w_116_116, w_060_125, w_075_087);
  or2  I116_137(w_116_137, w_053_004, w_008_067);
  and2 I116_191(w_116_191, w_025_013, w_104_303);
  nand2 I116_202(w_116_202, w_066_080, w_021_108);
  nand2 I116_208(w_116_208, w_084_122, w_028_042);
  and2 I116_214(w_116_214, w_114_278, w_059_445);
  nand2 I116_218(w_116_218, w_024_123, w_052_035);
  nand2 I116_243(w_116_243, w_043_026, w_047_368);
  or2  I116_275(w_116_275, w_018_288, w_108_008);
  nand2 I117_016(w_117_016, w_082_053, w_050_161);
  not1 I117_060(w_117_060, w_089_400);
  and2 I117_138(w_117_138, w_097_167, w_056_102);
  nand2 I117_157(w_117_157, w_071_235, w_010_334);
  not1 I117_161(w_117_161, w_027_086);
  and2 I117_176(w_117_176, w_015_002, w_052_086);
  nand2 I117_201(w_117_201, w_107_069, w_096_054);
  nand2 I117_221(w_117_221, w_104_223, w_110_142);
  nand2 I117_238(w_117_238, w_038_044, w_111_087);
  and2 I117_261(w_117_261, w_005_016, w_005_142);
  nand2 I117_266(w_117_266, w_110_161, w_069_028);
  or2  I117_279(w_117_279, w_059_121, w_092_123);
  not1 I117_289(w_117_289, w_109_000);
  not1 I117_294(w_117_294, w_051_132);
  or2  I117_322(w_117_322, w_074_003, w_115_320);
  not1 I117_324(w_117_324, w_088_030);
  and2 I117_325(w_117_325, w_063_013, w_062_004);
  and2 I117_341(w_117_341, w_086_001, w_113_075);
  nand2 I117_344(w_117_344, w_106_295, w_034_032);
  or2  I117_353(w_117_353, w_105_078, w_108_024);
  or2  I117_357(w_117_357, w_074_002, w_085_108);
  nand2 I117_362(w_117_362, w_086_038, w_114_022);
  or2  I117_375(w_117_375, w_049_320, w_098_013);
  not1 I117_386(w_117_386, w_007_084);
  nand2 I117_403(w_117_403, w_061_236, w_032_087);
  not1 I117_406(w_117_406, w_050_046);
  not1 I117_410(w_117_410, w_041_173);
  or2  I117_411(w_117_411, w_003_059, w_067_039);
  not1 I117_414(w_117_414, w_031_008);
  or2  I117_434(w_117_434, w_001_006, w_052_097);
  and2 I117_449(w_117_449, w_051_002, w_006_000);
  nand2 I118_020(w_118_020, w_060_220, w_066_131);
  or2  I118_024(w_118_024, w_066_113, w_039_225);
  not1 I118_026(w_118_026, w_025_097);
  and2 I118_046(w_118_046, w_009_056, w_081_084);
  nand2 I118_054(w_118_054, w_051_060, w_070_000);
  not1 I118_060(w_118_060, w_032_102);
  and2 I118_080(w_118_080, w_017_072, w_037_127);
  or2  I118_084(w_118_084, w_043_019, w_015_080);
  not1 I118_104(w_118_104, w_029_232);
  or2  I118_108(w_118_108, w_087_279, w_039_014);
  not1 I118_141(w_118_141, w_036_261);
  not1 I118_172(w_118_172, w_043_069);
  nand2 I118_175(w_118_175, w_061_072, w_096_146);
  or2  I118_187(w_118_187, w_061_208, w_112_184);
  or2  I118_194(w_118_194, w_053_026, w_044_023);
  or2  I118_196(w_118_196, w_034_129, w_065_007);
  nand2 I118_217(w_118_217, w_085_139, w_054_113);
  or2  I118_242(w_118_242, w_024_131, w_040_002);
  and2 I118_277(w_118_277, w_047_090, w_110_049);
  or2  I118_293(w_118_293, w_020_005, w_105_026);
  or2  I118_297(w_118_297, w_028_184, w_072_073);
  and2 I118_310(w_118_310, w_063_020, w_017_042);
  not1 I118_329(w_118_329, w_056_111);
  not1 I119_001(w_119_001, w_076_020);
  and2 I119_006(w_119_006, w_039_182, w_095_052);
  nand2 I119_040(w_119_040, w_031_045, w_093_281);
  and2 I119_101(w_119_101, w_028_345, w_068_066);
  not1 I119_107(w_119_107, w_026_098);
  not1 I119_114(w_119_114, w_105_012);
  or2  I119_122(w_119_122, w_004_182, w_068_042);
  and2 I119_136(w_119_136, w_113_042, w_014_022);
  or2  I119_141(w_119_141, w_013_154, w_038_093);
  not1 I119_157(w_119_157, w_011_251);
  or2  I119_168(w_119_168, w_065_159, w_116_214);
  not1 I119_184(w_119_184, w_076_062);
  nand2 I119_187(w_119_187, w_087_142, w_094_028);
  not1 I119_222(w_119_222, w_080_011);
  not1 I119_250(w_119_250, w_059_133);
  not1 I119_279(w_119_279, w_080_023);
  and2 I119_282(w_119_282, w_084_132, w_074_004);
  and2 I119_287(w_119_287, w_037_053, w_112_363);
  or2  I120_004(w_120_004, w_089_288, w_014_049);
  not1 I120_009(w_120_009, w_106_342);
  nand2 I120_016(w_120_016, w_082_101, w_031_011);
  not1 I120_021(w_120_021, w_097_139);
  nand2 I120_040(w_120_040, w_082_038, w_091_189);
  not1 I120_043(w_120_043, w_051_210);
  or2  I120_045(w_120_045, w_043_064, w_073_044);
  and2 I120_061(w_120_061, w_030_061, w_078_011);
  not1 I120_063(w_120_063, w_056_141);
  or2  I120_064(w_120_064, w_054_034, w_053_022);
  or2  I120_065(w_120_065, w_000_091, w_009_048);
  nand2 I120_070(w_120_070, w_040_005, w_055_048);
  or2  I120_086(w_120_086, w_049_272, w_038_037);
  not1 I120_088(w_120_088, w_025_146);
  or2  I120_089(w_120_089, w_050_058, w_090_068);
  nand2 I120_092(w_120_092, w_047_224, w_016_117);
  or2  I120_109(w_120_109, w_035_061, w_019_037);
  or2  I120_110(w_120_110, w_059_284, w_068_012);
  and2 I120_115(w_120_115, w_037_058, w_107_058);
  nand2 I120_117(w_120_117, w_047_278, w_077_024);
  not1 I120_136(w_120_136, w_085_017);
  and2 I120_140(w_120_140, w_078_006, w_072_096);
  nand2 I120_168(w_120_168, w_070_034, w_022_046);
  and2 I120_193(w_120_193, w_050_001, w_001_004);
  and2 I121_001(w_121_001, w_115_164, w_101_052);
  or2  I121_034(w_121_034, w_116_054, w_089_416);
  not1 I121_035(w_121_035, w_078_078);
  and2 I121_054(w_121_054, w_117_353, w_081_027);
  and2 I121_070(w_121_070, w_028_041, w_054_211);
  not1 I121_090(w_121_090, w_012_012);
  and2 I121_096(w_121_096, w_120_070, w_066_038);
  nand2 I121_107(w_121_107, w_106_164, w_117_266);
  not1 I121_126(w_121_126, w_018_026);
  nand2 I121_128(w_121_128, w_057_007, w_090_287);
  nand2 I121_159(w_121_159, w_018_125, w_056_110);
  not1 I121_164(w_121_164, w_017_029);
  or2  I121_242(w_121_242, w_099_110, w_118_104);
  nand2 I121_247(w_121_247, w_099_123, w_037_050);
  and2 I121_269(w_121_269, w_012_068, w_117_324);
  nand2 I121_284(w_121_284, w_042_145, w_051_016);
  nand2 I121_300(w_121_300, w_086_052, w_100_157);
  nand2 I122_002(w_122_002, w_024_042, w_112_108);
  nand2 I122_004(w_122_004, w_094_014, w_008_088);
  or2  I122_014(w_122_014, w_092_005, w_016_051);
  or2  I122_021(w_122_021, w_089_074, w_096_174);
  or2  I122_026(w_122_026, w_108_017, w_050_111);
  nand2 I122_028(w_122_028, w_017_059, w_097_027);
  nand2 I122_034(w_122_034, w_062_002, w_008_119);
  or2  I122_045(w_122_045, w_101_329, w_013_187);
  nand2 I122_057(w_122_057, w_009_058, w_026_334);
  and2 I122_079(w_122_079, w_031_007, w_042_033);
  not1 I122_084(w_122_084, w_091_123);
  not1 I122_086(w_122_086, w_109_000);
  not1 I122_089(w_122_089, w_029_098);
  nand2 I122_092(w_122_092, w_018_164, w_110_041);
  nand2 I122_096(w_122_096, w_035_084, w_002_020);
  or2  I122_107(w_122_107, w_034_238, w_118_196);
  not1 I122_110(w_122_110, w_034_066);
  or2  I122_113(w_122_113, w_086_042, w_074_004);
  not1 I122_114(w_122_114, w_070_047);
  or2  I122_125(w_122_125, w_098_005, w_022_116);
  not1 I122_128(w_122_128, w_013_073);
  and2 I122_141(w_122_141, w_027_201, w_022_139);
  not1 I122_152(w_122_152, w_116_026);
  and2 I122_157(w_122_157, w_058_025, w_067_004);
  not1 I122_161(w_122_161, w_081_029);
  not1 I122_163(w_122_163, w_108_050);
  or2  I123_007(w_123_007, w_103_001, w_020_176);
  and2 I123_012(w_123_012, w_057_005, w_097_070);
  and2 I123_023(w_123_023, w_041_109, w_068_025);
  nand2 I123_026(w_123_026, w_014_221, w_066_154);
  not1 I123_030(w_123_030, w_043_113);
  not1 I123_055(w_123_055, w_111_037);
  not1 I123_062(w_123_062, w_113_020);
  or2  I123_067(w_123_067, w_081_035, w_054_177);
  and2 I123_068(w_123_068, w_086_158, w_002_022);
  or2  I123_075(w_123_075, w_046_090, w_067_001);
  and2 I123_077(w_123_077, w_106_380, w_102_097);
  not1 I123_078(w_123_078, w_051_110);
  or2  I123_082(w_123_082, w_091_264, w_098_005);
  not1 I123_087(w_123_087, w_066_097);
  nand2 I123_120(w_123_120, w_041_160, w_046_182);
  and2 I123_124(w_123_124, w_010_005, w_030_062);
  or2  I123_149(w_123_149, w_087_314, w_048_366);
  and2 I123_167(w_123_167, w_009_025, w_085_065);
  nand2 I123_188(w_123_188, w_087_083, w_112_033);
  or2  I123_210(w_123_210, w_044_036, w_051_198);
  and2 I123_255(w_123_255, w_029_068, w_021_049);
  not1 I123_265(w_123_265, w_082_141);
  not1 I123_296(w_123_296, w_121_164);
  and2 I123_326(w_123_326, w_116_094, w_122_161);
  or2  I124_001(w_124_001, w_044_136, w_114_098);
  not1 I124_002(w_124_002, w_033_013);
  nand2 I124_020(w_124_020, w_107_046, w_083_179);
  nand2 I124_030(w_124_030, w_008_057, w_053_022);
  and2 I124_031(w_124_031, w_091_417, w_068_055);
  and2 I124_078(w_124_078, w_015_047, w_089_442);
  nand2 I124_088(w_124_088, w_060_049, w_091_411);
  not1 I124_099(w_124_099, w_066_135);
  not1 I124_106(w_124_106, w_021_009);
  nand2 I124_116(w_124_116, w_059_293, w_029_086);
  or2  I124_147(w_124_147, w_062_020, w_089_189);
  or2  I124_162(w_124_162, w_075_074, w_030_091);
  nand2 I124_174(w_124_174, w_115_195, w_078_163);
  and2 I124_211(w_124_211, w_028_313, w_089_096);
  nand2 I124_234(w_124_234, w_084_337, w_057_058);
  not1 I125_010(w_125_010, w_027_123);
  and2 I125_030(w_125_030, w_119_168, w_085_044);
  not1 I125_081(w_125_081, w_040_006);
  nand2 I125_117(w_125_117, w_054_125, w_079_158);
  nand2 I125_132(w_125_132, w_075_024, w_034_267);
  and2 I125_152(w_125_152, w_052_058, w_019_048);
  not1 I125_165(w_125_165, w_064_053);
  and2 I125_166(w_125_166, w_029_245, w_104_061);
  nand2 I125_186(w_125_186, w_071_004, w_032_195);
  and2 I125_222(w_125_222, w_090_019, w_007_166);
  or2  I125_234(w_125_234, w_070_068, w_067_033);
  nand2 I125_239(w_125_239, w_012_046, w_063_024);
  nand2 I125_246(w_125_246, w_039_107, w_046_108);
  nand2 I125_249(w_125_249, w_046_113, w_077_113);
  nand2 I125_255(w_125_255, w_014_154, w_031_015);
  or2  I125_359(w_125_359, w_074_001, w_085_098);
  not1 I125_396(w_125_396, w_123_030);
  not1 I125_411(w_125_411, w_103_009);
  and2 I125_463(w_125_463, w_089_243, w_056_170);
  or2  I126_001(w_126_001, w_029_077, w_076_013);
  nand2 I126_005(w_126_005, w_069_026, w_034_179);
  not1 I126_009(w_126_009, w_017_063);
  or2  I126_012(w_126_012, w_082_196, w_014_248);
  nand2 I126_016(w_126_016, w_096_184, w_005_145);
  not1 I126_020(w_126_020, w_021_016);
  and2 I126_024(w_126_024, w_016_310, w_008_280);
  nand2 I126_036(w_126_036, w_111_048, w_041_077);
  not1 I126_040(w_126_040, w_084_327);
  and2 I127_016(w_127_016, w_006_000, w_100_179);
  nand2 I127_021(w_127_021, w_126_024, w_063_122);
  or2  I127_033(w_127_033, w_114_092, w_032_027);
  and2 I127_075(w_127_075, w_057_041, w_007_001);
  not1 I127_133(w_127_133, w_068_090);
  nand2 I127_140(w_127_140, w_101_145, w_040_005);
  not1 I127_172(w_127_172, w_115_247);
  or2  I127_189(w_127_189, w_108_010, w_004_066);
  nand2 I127_237(w_127_237, w_072_074, w_064_060);
  not1 I127_246(w_127_246, w_112_053);
  nand2 I127_256(w_127_256, w_093_269, w_044_036);
  or2  I127_260(w_127_260, w_055_065, w_007_377);
  nand2 I127_272(w_127_272, w_004_061, w_003_025);
  not1 I127_328(w_127_328, w_123_265);
  nand2 I127_368(w_127_368, w_117_294, w_007_266);
  or2  I127_371(w_127_371, w_070_061, w_040_000);
  nand2 I127_404(w_127_404, w_075_041, w_068_150);
  not1 I127_491(w_127_493, w_127_492);
  not1 I127_492(w_127_494, w_127_493);
  or2  I127_493(w_127_495, w_127_494, w_059_260);
  not1 I127_494(w_127_496, w_127_495);
  nand2 I127_495(w_127_497, w_127_496, w_077_120);
  nand2 I127_496(w_127_498, w_127_497, w_070_065);
  not1 I127_497(w_127_499, w_127_498);
  or2  I127_498(w_127_500, w_127_499, w_016_210);
  nand2 I127_499(w_127_501, w_127_500, w_033_027);
  not1 I127_500(w_127_502, w_127_501);
  or2  I127_501(w_127_503, w_127_502, w_064_053);
  and2 I127_502(w_127_492, w_127_503, w_115_212);
  and2 I127_503(w_127_508, w_039_056, w_127_507);
  or2  I127_504(w_127_509, w_065_035, w_127_508);
  not1 I127_505(w_127_510, w_127_509);
  and2 I127_506(w_127_511, w_043_043, w_127_510);
  nand2 I127_507(w_127_512, w_070_024, w_127_511);
  or2  I127_508(w_127_513, w_106_079, w_127_512);
  not1 I127_509(w_127_514, w_127_513);
  nand2 I127_510(w_127_515, w_127_534, w_127_514);
  nand2 I127_511(w_127_516, w_002_001, w_127_515);
  or2  I127_512(w_127_517, w_127_516, w_066_072);
  or2  I127_513(w_127_507, w_127_517, w_022_041);
  or2  I127_514(w_127_522, w_127_521, w_017_190);
  or2  I127_515(w_127_523, w_127_522, w_078_071);
  nand2 I127_516(w_127_524, w_127_523, w_074_002);
  nand2 I127_517(w_127_525, w_127_524, w_077_174);
  or2  I127_518(w_127_526, w_075_025, w_127_525);
  and2 I127_519(w_127_527, w_021_037, w_127_526);
  or2  I127_520(w_127_528, w_055_002, w_127_527);
  not1 I127_521(w_127_529, w_127_528);
  not1 I127_522(w_127_530, w_127_529);
  and2 I127_523(w_127_531, w_118_020, w_127_530);
  or2  I127_524(w_127_532, w_127_531, w_036_098);
  not1 I127_525(w_127_521, w_127_515);
  and2 I127_526(w_127_534, w_121_096, w_127_532);
  not1 I128_013(w_128_013, w_098_023);
  not1 I128_015(w_128_015, w_124_162);
  not1 I128_025(w_128_025, w_003_043);
  not1 I128_031(w_128_031, w_006_000);
  or2  I128_032(w_128_032, w_088_270, w_052_022);
  not1 I128_034(w_128_034, w_008_196);
  and2 I128_038(w_128_038, w_061_242, w_101_175);
  or2  I128_042(w_128_042, w_099_159, w_081_039);
  or2  I128_043(w_128_043, w_089_092, w_100_180);
  and2 I128_045(w_128_045, w_049_149, w_056_043);
  or2  I128_048(w_128_048, w_075_020, w_054_018);
  and2 I128_051(w_128_051, w_055_029, w_080_020);
  not1 I128_054(w_128_054, w_059_100);
  not1 I128_057(w_128_057, w_122_089);
  nand2 I128_058(w_128_058, w_008_064, w_095_080);
  and2 I128_061(w_127_505, w_125_010, w_127_492);
  and2 I128_062(w_127_519, w_127_505, w_127_507);
  not1 I129_000(w_129_000, w_127_519);
  not1 I130_009(w_130_009, w_002_012);
  not1 I130_012(w_130_012, w_067_000);
  or2  I130_021(w_130_021, w_083_002, w_008_017);
  nand2 I130_027(w_130_027, w_120_092, w_014_178);
  or2  I130_034(w_130_034, w_019_047, w_077_085);
  nand2 I130_037(w_130_037, w_067_004, w_019_027);
  and2 I130_068(w_130_068, w_103_018, w_104_260);
  or2  I130_072(w_130_072, w_100_312, w_087_067);
  or2  I130_086(w_130_086, w_099_038, w_053_021);
  and2 I130_087(w_130_087, w_021_041, w_041_135);
  nand2 I130_106(w_130_106, w_116_191, w_122_084);
  not1 I130_107(w_130_107, w_049_070);
  and2 I130_111(w_130_111, w_098_016, w_044_302);
  nand2 I130_137(w_130_137, w_081_020, w_122_014);
  not1 I130_142(w_130_142, w_059_280);
  nand2 I130_146(w_130_146, w_102_147, w_044_055);
  and2 I130_171(w_130_171, w_116_059, w_104_031);
  or2  I131_001(w_131_001, w_000_254, w_080_011);
  not1 I131_009(w_131_009, w_112_071);
  not1 I131_012(w_131_012, w_015_050);
  not1 I131_024(w_131_024, w_020_020);
  and2 I131_040(w_131_040, w_051_046, w_013_040);
  nand2 I131_041(w_131_041, w_077_135, w_057_036);
  nand2 I131_058(w_131_058, w_114_001, w_020_085);
  nand2 I131_063(w_131_063, w_108_030, w_099_180);
  nand2 I131_081(w_131_081, w_130_086, w_127_256);
  not1 I131_127(w_131_127, w_080_035);
  and2 I131_141(w_131_141, w_068_051, w_039_396);
  not1 I131_142(w_131_142, w_082_027);
  not1 I131_169(w_131_169, w_047_022);
  nand2 I131_191(w_131_191, w_009_203, w_086_195);
  or2  I131_196(w_131_196, w_115_203, w_038_008);
  or2  I131_198(w_131_198, w_000_431, w_072_042);
  not1 I132_037(w_132_037, w_123_255);
  and2 I132_054(w_132_054, w_049_079, w_110_051);
  nand2 I132_067(w_132_067, w_114_058, w_107_010);
  nand2 I132_100(w_132_100, w_114_195, w_072_075);
  nand2 I132_104(w_132_104, w_005_017, w_059_056);
  and2 I132_113(w_132_113, w_114_027, w_123_326);
  not1 I132_114(w_132_114, w_014_211);
  nand2 I132_133(w_132_133, w_074_003, w_112_073);
  or2  I132_169(w_132_169, w_125_222, w_063_030);
  or2  I132_176(w_132_176, w_055_018, w_074_000);
  nand2 I132_182(w_132_182, w_090_194, w_048_132);
  or2  I132_185(w_132_185, w_126_009, w_115_037);
  or2  I133_026(w_133_026, w_031_021, w_000_434);
  nand2 I133_068(w_133_068, w_041_096, w_079_193);
  and2 I133_076(w_133_076, w_102_078, w_037_018);
  nand2 I133_101(w_133_101, w_026_345, w_094_081);
  or2  I133_174(w_133_174, w_068_136, w_041_140);
  not1 I133_227(w_133_227, w_082_005);
  and2 I133_232(w_133_232, w_028_128, w_063_226);
  nand2 I133_282(w_133_282, w_092_065, w_052_056);
  nand2 I133_357(w_133_357, w_008_004, w_068_100);
  or2  I134_002(w_134_002, w_108_011, w_093_276);
  nand2 I134_003(w_134_003, w_074_005, w_127_075);
  and2 I134_004(w_134_004, w_040_002, w_003_086);
  not1 I134_020(w_134_020, w_111_066);
  not1 I134_022(w_134_022, w_047_259);
  not1 I134_026(w_134_026, w_122_057);
  or2  I134_033(w_134_033, w_038_077, w_042_001);
  not1 I134_034(w_134_034, w_061_094);
  not1 I134_042(w_134_042, w_119_250);
  and2 I134_043(w_134_043, w_105_167, w_059_004);
  nand2 I134_046(w_134_046, w_039_475, w_084_037);
  and2 I134_047(w_134_047, w_129_000, w_010_333);
  not1 I134_053(w_134_053, w_006_000);
  not1 I134_054(w_134_054, w_024_002);
  or2  I134_062(w_134_062, w_123_007, w_050_026);
  or2  I134_063(w_134_063, w_130_111, w_071_270);
  nand2 I134_064(w_134_064, w_044_163, w_094_155);
  not1 I134_068(w_134_068, w_029_133);
  nand2 I134_069(w_134_069, w_067_062, w_060_142);
  not1 I134_073(w_134_073, w_078_041);
  not1 I134_075(w_134_075, w_100_298);
  not1 I134_085(w_134_085, w_016_234);
  and2 I135_027(w_135_027, w_051_159, w_054_178);
  and2 I135_049(w_135_049, w_114_181, w_042_154);
  and2 I135_097(w_135_097, w_083_004, w_057_001);
  not1 I135_113(w_135_113, w_024_183);
  nand2 I135_115(w_135_115, w_101_158, w_083_090);
  nand2 I135_123(w_135_123, w_077_184, w_091_225);
  nand2 I135_131(w_135_131, w_046_086, w_092_109);
  or2  I135_153(w_135_153, w_123_023, w_075_054);
  nand2 I135_186(w_135_186, w_016_094, w_073_125);
  not1 I135_203(w_135_203, w_130_009);
  not1 I135_222(w_135_222, w_105_001);
  nand2 I135_250(w_135_250, w_021_070, w_035_096);
  and2 I136_001(w_136_001, w_048_079, w_118_172);
  nand2 I136_002(w_136_002, w_067_015, w_036_219);
  and2 I136_007(w_136_007, w_135_131, w_051_238);
  or2  I136_013(w_136_013, w_076_021, w_093_143);
  not1 I136_014(w_136_014, w_008_233);
  or2  I136_017(w_136_017, w_055_000, w_050_063);
  not1 I136_018(w_136_018, w_011_086);
  not1 I136_019(w_136_019, w_103_008);
  and2 I136_021(w_136_021, w_094_023, w_121_300);
  and2 I136_022(w_136_022, w_099_226, w_082_188);
  not1 I136_029(w_136_029, w_052_006);
  and2 I137_008(w_137_008, w_057_031, w_131_012);
  and2 I137_010(w_137_010, w_026_212, w_054_029);
  and2 I137_014(w_137_014, w_081_025, w_070_074);
  nand2 I137_021(w_137_021, w_042_200, w_023_156);
  and2 I137_031(w_137_031, w_113_066, w_022_091);
  and2 I137_035(w_137_035, w_135_097, w_056_176);
  not1 I137_041(w_137_041, w_102_003);
  and2 I137_045(w_137_045, w_086_102, w_015_068);
  or2  I137_050(w_137_050, w_047_185, w_102_044);
  and2 I137_054(w_137_054, w_080_015, w_121_035);
  and2 I137_057(w_137_057, w_126_001, w_020_007);
  nand2 I138_006(w_138_006, w_043_032, w_064_024);
  nand2 I138_013(w_138_013, w_065_133, w_075_130);
  nand2 I138_122(w_138_122, w_045_125, w_103_008);
  or2  I138_128(w_138_128, w_007_137, w_113_039);
  nand2 I138_174(w_138_174, w_094_357, w_088_397);
  and2 I138_215(w_138_215, w_098_008, w_114_050);
  or2  I138_217(w_138_217, w_027_057, w_004_314);
  and2 I138_223(w_138_223, w_060_060, w_005_115);
  and2 I138_240(w_138_242, w_138_241, w_048_143);
  or2  I138_241(w_138_243, w_071_191, w_138_242);
  and2 I138_242(w_138_244, w_138_259, w_138_243);
  nand2 I138_243(w_138_245, w_138_244, w_050_187);
  nand2 I138_244(w_138_246, w_138_245, w_136_002);
  not1 I138_245(w_138_247, w_138_246);
  not1 I138_246(w_138_248, w_138_247);
  not1 I138_247(w_138_241, w_138_248);
  nand2 I138_248(w_138_253, w_138_252, w_083_084);
  or2  I138_249(w_138_254, w_129_000, w_138_253);
  and2 I138_250(w_138_255, w_054_191, w_138_254);
  nand2 I138_251(w_138_256, w_138_255, w_102_076);
  or2  I138_252(w_138_257, w_138_256, w_014_058);
  not1 I138_253(w_138_252, w_138_244);
  and2 I138_254(w_138_259, w_002_013, w_138_257);
  and2 I139_016(w_139_016, w_107_069, w_050_042);
  or2  I139_025(w_139_025, w_103_006, w_026_018);
  or2  I139_030(w_139_030, w_134_033, w_082_134);
  nand2 I139_043(w_139_043, w_004_142, w_099_054);
  or2  I139_112(w_139_112, w_001_003, w_031_038);
  or2  I139_150(w_139_150, w_101_305, w_001_006);
  and2 I139_154(w_139_154, w_050_026, w_051_056);
  not1 I139_164(w_139_164, w_009_015);
  and2 I139_176(w_139_176, w_009_001, w_061_284);
  nand2 I139_182(w_139_182, w_038_031, w_030_045);
  and2 I139_187(w_139_187, w_120_086, w_125_165);
  nand2 I139_188(w_139_188, w_012_265, w_100_194);
  nand2 I139_228(w_139_230, w_044_133, w_139_229);
  or2  I139_229(w_139_231, w_112_232, w_139_230);
  and2 I139_230(w_139_229, w_070_095, w_139_231);
  nand2 I140_005(w_140_005, w_054_165, w_033_037);
  not1 I140_026(w_140_026, w_091_235);
  not1 I140_043(w_140_043, w_058_037);
  nand2 I140_044(w_140_044, w_087_178, w_096_030);
  and2 I140_049(w_140_049, w_118_060, w_089_380);
  nand2 I140_071(w_140_071, w_115_242, w_131_012);
  and2 I140_080(w_140_080, w_117_221, w_113_042);
  not1 I140_084(w_140_084, w_105_035);
  nand2 I140_106(w_140_106, w_136_001, w_051_266);
  or2  I140_110(w_140_110, w_091_289, w_054_090);
  nand2 I140_157(w_140_157, w_113_059, w_112_017);
  or2  I140_196(w_140_196, w_087_217, w_131_001);
  nand2 I140_266(w_140_266, w_003_089, w_059_390);
  not1 I140_300(w_140_300, w_096_022);
  nand2 I141_005(w_141_005, w_070_065, w_132_114);
  not1 I141_022(w_141_022, w_074_004);
  or2  I141_061(w_141_061, w_044_295, w_077_029);
  nand2 I141_122(w_141_122, w_072_022, w_087_147);
  and2 I141_153(w_141_153, w_033_051, w_003_094);
  and2 I141_154(w_141_154, w_099_015, w_086_068);
  not1 I141_163(w_141_163, w_081_030);
  or2  I141_169(w_141_169, w_022_016, w_109_001);
  not1 I141_172(w_141_172, w_107_069);
  not1 I141_193(w_141_193, w_071_010);
  nand2 I141_207(w_141_207, w_079_452, w_028_032);
  not1 I141_261(w_141_261, w_097_205);
  and2 I142_000(w_142_000, w_117_161, w_061_050);
  and2 I142_070(w_142_070, w_132_169, w_136_014);
  or2  I142_078(w_142_078, w_057_048, w_011_059);
  not1 I142_083(w_142_083, w_094_033);
  not1 I142_086(w_142_086, w_114_038);
  not1 I142_098(w_142_098, w_070_009);
  or2  I142_103(w_142_103, w_061_178, w_073_040);
  not1 I142_106(w_142_106, w_097_146);
  nand2 I142_111(w_142_111, w_118_194, w_111_020);
  nand2 I142_116(w_142_116, w_007_018, w_117_157);
  nand2 I142_122(w_142_122, w_043_238, w_119_114);
  nand2 I142_131(w_142_131, w_056_147, w_093_351);
  not1 I142_146(w_142_146, w_132_182);
  not1 I142_150(w_142_150, w_009_005);
  or2  I142_173(w_142_173, w_037_086, w_127_237);
  nand2 I142_176(w_142_176, w_041_036, w_006_000);
  nand2 I142_204(w_142_204, w_049_182, w_052_047);
  not1 I142_250(w_142_250, w_128_015);
  and2 I142_279(w_142_279, w_111_048, w_127_328);
  not1 I142_303(w_142_303, w_106_408);
  not1 I143_002(w_143_002, w_104_365);
  not1 I143_018(w_143_018, w_031_063);
  or2  I143_025(w_143_025, w_046_210, w_121_090);
  or2  I143_033(w_143_033, w_136_001, w_021_098);
  or2  I143_054(w_143_054, w_104_192, w_107_021);
  and2 I143_061(w_143_061, w_134_064, w_031_025);
  or2  I143_070(w_143_070, w_054_056, w_064_046);
  and2 I143_087(w_143_087, w_057_051, w_080_005);
  not1 I143_088(w_143_088, w_000_448);
  or2  I143_092(w_143_092, w_101_034, w_013_024);
  nand2 I143_099(w_143_099, w_040_002, w_026_058);
  and2 I143_103(w_143_103, w_125_132, w_041_271);
  nand2 I143_107(w_143_107, w_004_130, w_132_037);
  and2 I144_004(w_144_004, w_131_009, w_110_027);
  or2  I144_010(w_144_010, w_101_099, w_093_269);
  or2  I144_016(w_144_016, w_118_084, w_130_107);
  not1 I144_045(w_144_045, w_032_137);
  and2 I144_058(w_144_058, w_092_076, w_140_071);
  and2 I144_062(w_144_062, w_059_262, w_129_000);
  and2 I144_064(w_144_064, w_109_000, w_013_060);
  nand2 I144_095(w_144_095, w_078_055, w_024_169);
  or2  I144_105(w_144_105, w_008_092, w_128_048);
  not1 I144_107(w_144_107, w_129_000);
  or2  I144_124(w_144_124, w_126_040, w_111_055);
  nand2 I144_136(w_144_136, w_021_106, w_004_190);
  or2  I144_151(w_144_151, w_093_272, w_083_031);
  or2  I144_172(w_144_172, w_128_057, w_002_005);
  and2 I144_186(w_144_186, w_059_297, w_001_003);
  not1 I145_006(w_145_006, w_084_076);
  nand2 I145_009(w_145_009, w_080_013, w_087_074);
  not1 I145_063(w_145_063, w_128_045);
  nand2 I145_072(w_145_072, w_099_052, w_064_058);
  nand2 I145_073(w_145_073, w_113_002, w_011_222);
  not1 I145_143(w_145_143, w_016_253);
  or2  I145_196(w_145_196, w_137_057, w_142_250);
  not1 I145_215(w_145_215, w_137_054);
  or2  I145_219(w_145_219, w_012_218, w_084_176);
  nand2 I145_250(w_145_250, w_141_172, w_123_296);
  nand2 I145_333(w_145_333, w_083_023, w_124_234);
  and2 I145_393(w_145_393, w_015_027, w_029_179);
  and2 I146_011(w_146_011, w_060_379, w_135_222);
  not1 I146_017(w_146_017, w_000_376);
  and2 I146_033(w_146_033, w_017_138, w_112_050);
  not1 I146_037(w_146_037, w_102_013);
  nand2 I146_041(w_146_041, w_044_172, w_104_379);
  and2 I146_050(w_146_050, w_051_042, w_144_172);
  or2  I146_061(w_146_061, w_122_079, w_026_103);
  or2  I146_064(w_146_064, w_032_000, w_086_120);
  and2 I146_087(w_146_087, w_101_106, w_097_064);
  and2 I146_161(w_146_161, w_050_070, w_026_022);
  or2  I146_168(w_146_168, w_100_003, w_044_087);
  not1 I146_200(w_146_200, w_090_298);
  nand2 I146_220(w_146_220, w_096_030, w_087_148);
  not1 I146_228(w_146_228, w_126_005);
  nand2 I146_245(w_146_245, w_074_003, w_117_386);
  or2  I146_307(w_146_307, w_119_279, w_099_075);
  or2  I147_012(w_147_012, w_011_135, w_044_133);
  not1 I147_019(w_147_019, w_119_136);
  or2  I147_033(w_147_033, w_114_077, w_017_030);
  and2 I147_063(w_147_063, w_120_193, w_112_304);
  and2 I147_066(w_147_066, w_024_073, w_048_072);
  or2  I147_074(w_147_074, w_056_163, w_104_327);
  not1 I147_084(w_147_084, w_012_135);
  and2 I147_106(w_147_106, w_087_082, w_127_016);
  and2 I147_107(w_147_107, w_124_030, w_038_099);
  nand2 I147_119(w_147_119, w_012_098, w_141_169);
  and2 I147_127(w_147_127, w_005_191, w_026_209);
  nand2 I147_129(w_147_129, w_039_364, w_084_111);
  not1 I147_136(w_147_136, w_108_046);
  not1 I147_138(w_147_138, w_120_089);
  or2  I147_151(w_147_151, w_015_020, w_138_174);
  and2 I147_175(w_147_175, w_077_246, w_118_026);
  not1 I147_191(w_147_191, w_001_004);
  not1 I148_012(w_148_012, w_010_025);
  not1 I148_022(w_148_022, w_085_079);
  or2  I148_028(w_148_028, w_114_057, w_034_146);
  or2  I148_038(w_148_038, w_090_111, w_129_000);
  not1 I148_069(w_148_069, w_009_139);
  or2  I148_073(w_148_073, w_118_020, w_037_086);
  not1 I148_087(w_148_087, w_091_070);
  not1 I148_121(w_148_121, w_000_005);
  and2 I148_129(w_148_129, w_012_349, w_024_151);
  and2 I148_242(w_148_242, w_021_011, w_032_074);
  or2  I148_251(w_148_251, w_120_065, w_050_188);
  and2 I148_324(w_148_324, w_113_048, w_118_277);
  and2 I149_000(w_149_000, w_002_024, w_090_281);
  nand2 I149_001(w_149_001, w_093_107, w_099_022);
  and2 I149_003(w_149_003, w_015_067, w_134_073);
  and2 I149_004(w_149_004, w_102_155, w_087_138);
  nand2 I149_005(w_149_005, w_001_005, w_071_352);
  or2  I149_007(w_149_007, w_146_307, w_044_154);
  or2  I149_008(w_149_008, w_084_286, w_010_251);
  not1 I149_011(w_149_011, w_002_019);
  not1 I149_018(w_149_018, w_136_013);
  or2  I149_019(w_149_019, w_108_010, w_082_221);
  nand2 I149_022(w_149_022, w_026_232, w_068_014);
  nand2 I149_023(w_149_023, w_144_095, w_018_322);
  and2 I149_024(w_149_024, w_072_067, w_007_073);
  not1 I149_026(w_149_026, w_001_000);
  and2 I149_027(w_149_027, w_052_056, w_061_383);
  and2 I149_028(w_149_028, w_037_069, w_090_288);
  and2 I150_024(w_150_024, w_137_031, w_068_040);
  and2 I150_063(w_150_063, w_128_051, w_102_071);
  and2 I150_082(w_150_082, w_003_096, w_041_288);
  and2 I150_089(w_150_089, w_061_014, w_076_011);
  or2  I150_106(w_150_106, w_061_406, w_059_072);
  or2  I150_122(w_150_122, w_146_220, w_024_000);
  or2  I150_146(w_150_146, w_120_064, w_123_077);
  nand2 I150_156(w_150_156, w_101_249, w_120_063);
  or2  I150_176(w_150_176, w_116_022, w_129_000);
  and2 I150_225(w_150_225, w_032_006, w_052_013);
  or2  I150_320(w_150_320, w_059_359, w_124_001);
  or2  I150_334(w_150_334, w_043_119, w_007_240);
  or2  I150_392(w_150_392, w_022_126, w_030_089);
  not1 I151_000(w_151_000, w_086_165);
  or2  I151_007(w_151_007, w_059_041, w_142_204);
  nand2 I151_008(w_151_008, w_117_357, w_023_367);
  or2  I151_010(w_151_010, w_076_062, w_117_176);
  not1 I151_021(w_151_021, w_104_301);
  nand2 I151_023(w_151_023, w_061_174, w_075_089);
  nand2 I151_029(w_151_029, w_040_004, w_084_214);
  not1 I151_033(w_151_033, w_030_087);
  and2 I151_034(w_151_034, w_129_000, w_031_024);
  or2  I151_036(w_151_036, w_070_084, w_133_101);
  or2  I151_038(w_151_038, w_114_038, w_002_002);
  nand2 I151_041(w_151_041, w_031_002, w_069_031);
  and2 I152_022(w_152_022, w_077_236, w_144_058);
  or2  I152_029(w_152_029, w_109_000, w_018_130);
  and2 I152_032(w_152_032, w_096_165, w_117_449);
  or2  I152_050(w_152_050, w_118_024, w_031_011);
  or2  I152_053(w_152_053, w_090_111, w_126_005);
  or2  I152_056(w_152_056, w_106_022, w_114_115);
  or2  I152_059(w_152_059, w_102_083, w_111_007);
  not1 I152_062(w_152_062, w_096_296);
  and2 I152_072(w_152_072, w_084_113, w_006_000);
  nand2 I152_083(w_152_083, w_007_347, w_060_023);
  or2  I152_120(w_152_120, w_040_001, w_057_011);
  nand2 I152_132(w_152_132, w_147_119, w_007_041);
  and2 I152_134(w_152_134, w_040_002, w_107_022);
  or2  I152_147(w_152_147, w_125_411, w_029_073);
  and2 I152_191(w_152_191, w_028_000, w_144_105);
  and2 I153_001(w_153_001, w_131_040, w_090_262);
  nand2 I153_007(w_153_007, w_121_128, w_143_087);
  nand2 I153_008(w_153_008, w_106_422, w_097_008);
  and2 I153_025(w_153_025, w_009_019, w_054_199);
  and2 I153_093(w_153_093, w_092_176, w_117_325);
  not1 I153_108(w_153_108, w_000_012);
  and2 I153_125(w_153_125, w_141_022, w_062_006);
  not1 I153_186(w_153_186, w_009_149);
  not1 I153_209(w_153_209, w_009_121);
  and2 I153_218(w_153_218, w_069_091, w_015_060);
  and2 I153_255(w_153_255, w_149_008, w_150_024);
  and2 I153_297(w_153_297, w_138_006, w_014_132);
  not1 I153_331(w_153_331, w_019_048);
  not1 I153_409(w_153_409, w_110_210);
  or2  I153_424(w_153_424, w_147_033, w_091_168);
  or2  I153_461(w_153_461, w_001_005, w_078_032);
  and2 I154_009(w_154_009, w_098_006, w_001_006);
  not1 I154_013(w_154_013, w_098_013);
  nand2 I154_024(w_154_024, w_050_126, w_024_182);
  not1 I154_047(w_154_047, w_063_047);
  not1 I154_050(w_154_050, w_070_053);
  or2  I154_051(w_154_051, w_132_100, w_112_103);
  or2  I154_058(w_154_058, w_010_014, w_032_132);
  or2  I154_062(w_154_062, w_085_206, w_102_039);
  or2  I154_075(w_154_075, w_112_212, w_140_157);
  or2  I154_078(w_154_078, w_134_063, w_097_148);
  or2  I154_103(w_154_103, w_086_047, w_147_175);
  not1 I154_106(w_154_106, w_036_028);
  or2  I155_023(w_155_023, w_078_144, w_122_028);
  or2  I155_072(w_155_072, w_084_030, w_071_055);
  and2 I155_080(w_155_080, w_141_261, w_118_310);
  not1 I155_101(w_155_101, w_017_156);
  or2  I155_102(w_155_102, w_075_093, w_141_122);
  or2  I155_110(w_155_110, w_116_202, w_056_078);
  and2 I155_165(w_155_165, w_033_053, w_150_063);
  and2 I155_189(w_155_189, w_003_045, w_011_155);
  not1 I155_231(w_155_231, w_002_003);
  nand2 I155_237(w_155_237, w_098_015, w_043_171);
  and2 I155_261(w_155_261, w_019_013, w_143_002);
  not1 I155_272(w_155_272, w_088_335);
  nand2 I155_322(w_155_322, w_034_080, w_146_228);
  not1 I155_329(w_155_329, w_049_189);
  and2 I156_066(w_156_066, w_048_317, w_072_048);
  not1 I156_090(w_156_090, w_107_045);
  nand2 I156_115(w_156_115, w_152_050, w_065_027);
  and2 I156_144(w_156_144, w_103_018, w_068_119);
  and2 I156_153(w_156_153, w_118_297, w_101_163);
  and2 I156_168(w_156_168, w_095_030, w_102_028);
  and2 I156_217(w_156_217, w_096_039, w_044_034);
  nand2 I156_225(w_156_225, w_077_104, w_124_020);
  or2  I156_302(w_156_302, w_022_160, w_135_186);
  and2 I157_019(w_157_019, w_022_102, w_098_017);
  not1 I157_165(w_157_165, w_130_027);
  nand2 I157_229(w_157_229, w_035_101, w_014_259);
  and2 I157_242(w_157_242, w_010_364, w_089_032);
  and2 I157_393(w_157_393, w_070_017, w_118_187);
  not1 I157_434(w_157_434, w_097_133);
  and2 I158_000(w_158_000, w_143_088, w_103_005);
  not1 I158_001(w_158_001, w_005_186);
  not1 I158_003(w_158_003, w_144_045);
  or2  I158_006(w_158_006, w_032_073, w_023_047);
  and2 I158_007(w_158_007, w_036_078, w_085_197);
  and2 I158_011(w_158_011, w_123_087, w_035_109);
  and2 I158_013(w_158_013, w_027_086, w_006_000);
  nand2 I158_016(w_158_016, w_139_154, w_109_000);
  or2  I158_025(w_158_025, w_094_147, w_105_077);
  nand2 I158_027(w_158_027, w_090_317, w_096_134);
  not1 I158_036(w_158_036, w_002_011);
  or2  I158_037(w_158_039, w_005_219, w_158_038);
  nand2 I158_038(w_158_040, w_158_039, w_074_004);
  not1 I158_039(w_158_041, w_158_040);
  and2 I158_040(w_158_042, w_158_041, w_147_127);
  nand2 I158_041(w_158_043, w_158_042, w_101_039);
  nand2 I158_042(w_158_044, w_158_043, w_075_124);
  or2  I158_043(w_158_045, w_129_000, w_158_044);
  and2 I158_044(w_158_046, w_158_045, w_127_260);
  and2 I158_045(w_158_047, w_158_046, w_006_000);
  not1 I158_046(w_158_048, w_158_047);
  or2  I158_047(w_158_038, w_057_036, w_158_048);
  or2  I159_005(w_159_005, w_065_024, w_090_190);
  and2 I159_007(w_159_007, w_042_121, w_063_200);
  and2 I159_055(w_159_055, w_121_284, w_142_103);
  nand2 I159_072(w_159_072, w_067_023, w_118_217);
  not1 I159_073(w_159_073, w_149_008);
  not1 I159_080(w_159_080, w_081_061);
  and2 I159_092(w_159_092, w_014_114, w_114_208);
  or2  I159_107(w_159_107, w_156_144, w_030_178);
  or2  I159_128(w_159_128, w_049_060, w_112_081);
  nand2 I159_158(w_159_158, w_039_215, w_130_137);
  nand2 I159_199(w_159_199, w_021_024, w_057_050);
  not1 I159_210(w_159_210, w_058_020);
  and2 I160_013(w_160_013, w_159_080, w_014_017);
  nand2 I160_014(w_160_014, w_115_379, w_041_228);
  and2 I160_025(w_160_025, w_155_023, w_062_020);
  nand2 I160_060(w_160_060, w_104_007, w_143_033);
  or2  I160_071(w_160_071, w_069_144, w_145_333);
  or2  I160_072(w_160_072, w_143_025, w_129_000);
  or2  I160_075(w_160_075, w_117_414, w_111_015);
  nand2 I160_102(w_160_102, w_095_000, w_122_107);
  and2 I160_114(w_160_114, w_008_100, w_086_073);
  nand2 I160_132(w_160_132, w_011_231, w_142_279);
  and2 I160_138(w_160_138, w_134_068, w_115_032);
  and2 I161_013(w_161_013, w_037_069, w_082_088);
  and2 I161_031(w_161_031, w_044_050, w_010_256);
  not1 I161_039(w_161_039, w_131_198);
  not1 I161_067(w_161_067, w_010_042);
  or2  I161_083(w_161_083, w_084_062, w_085_002);
  nand2 I161_141(w_161_141, w_038_066, w_041_098);
  and2 I161_153(w_161_153, w_103_018, w_096_145);
  nand2 I161_160(w_161_160, w_108_019, w_086_024);
  and2 I161_171(w_161_171, w_063_222, w_124_099);
  and2 I161_207(w_161_207, w_082_103, w_082_125);
  nand2 I161_219(w_161_219, w_160_071, w_030_035);
  nand2 I161_261(w_161_261, w_065_072, w_018_089);
  not1 I162_000(w_162_000, w_134_003);
  not1 I162_001(w_162_001, w_012_045);
  nand2 I162_005(w_162_005, w_004_332, w_069_017);
  nand2 I162_007(w_162_007, w_106_482, w_060_011);
  nand2 I162_008(w_162_008, w_103_003, w_020_105);
  not1 I162_009(w_162_009, w_147_129);
  and2 I162_010(w_162_010, w_123_167, w_045_036);
  and2 I162_011(w_162_011, w_051_010, w_089_007);
  and2 I162_012(w_162_012, w_012_024, w_141_153);
  or2  I162_013(w_162_013, w_096_009, w_099_006);
  nand2 I162_014(w_162_014, w_013_194, w_092_016);
  not1 I162_015(w_162_015, w_128_042);
  nand2 I162_017(w_162_017, w_081_008, w_153_008);
  or2  I163_000(w_163_000, w_123_055, w_024_042);
  or2  I163_003(w_163_003, w_081_073, w_092_026);
  not1 I163_007(w_163_007, w_069_106);
  not1 I163_016(w_163_016, w_007_071);
  and2 I163_035(w_163_035, w_134_020, w_048_083);
  nand2 I163_054(w_163_054, w_142_122, w_000_033);
  and2 I163_070(w_163_070, w_083_056, w_005_125);
  or2  I163_133(w_163_133, w_073_101, w_116_191);
  not1 I163_147(w_163_147, w_001_005);
  nand2 I163_156(w_163_156, w_009_007, w_006_000);
  and2 I163_171(w_163_171, w_076_026, w_092_032);
  and2 I163_187(w_163_187, w_048_193, w_065_104);
  nand2 I163_210(w_163_210, w_024_114, w_009_040);
  and2 I163_250(w_163_250, w_091_258, w_021_092);
  and2 I163_330(w_163_330, w_129_000, w_016_113);
  not1 I163_371(w_163_371, w_105_121);
  not1 I163_383(w_163_383, w_059_264);
  nand2 I164_001(w_164_001, w_051_042, w_148_073);
  or2  I164_012(w_164_012, w_003_088, w_036_045);
  or2  I164_020(w_164_020, w_102_059, w_063_223);
  and2 I164_027(w_164_027, w_051_266, w_058_075);
  or2  I164_058(w_164_058, w_079_247, w_161_067);
  or2  I164_090(w_164_090, w_102_129, w_006_000);
  nand2 I164_098(w_164_098, w_101_105, w_134_062);
  and2 I164_106(w_164_106, w_003_008, w_083_079);
  nand2 I164_119(w_164_119, w_123_082, w_117_016);
  not1 I164_132(w_164_132, w_103_015);
  or2  I164_136(w_164_136, w_024_132, w_161_083);
  or2  I164_163(w_164_163, w_121_107, w_105_293);
  not1 I164_187(w_164_189, w_164_188);
  not1 I164_188(w_164_190, w_164_189);
  nand2 I164_189(w_164_191, w_139_150, w_164_190);
  not1 I164_190(w_164_192, w_164_191);
  or2  I164_191(w_164_193, w_084_270, w_164_192);
  nand2 I164_192(w_164_194, w_106_269, w_164_193);
  or2  I164_193(w_164_195, w_164_194, w_067_044);
  nand2 I164_194(w_164_188, w_164_195, w_051_172);
  nand2 I165_004(w_165_004, w_001_005, w_019_046);
  nand2 I165_028(w_165_028, w_100_062, w_161_039);
  not1 I165_057(w_165_057, w_127_140);
  nand2 I165_092(w_165_092, w_066_006, w_096_235);
  nand2 I165_104(w_165_104, w_004_057, w_118_080);
  and2 I165_111(w_165_111, w_042_196, w_025_244);
  and2 I165_112(w_165_112, w_147_138, w_139_112);
  or2  I165_174(w_165_174, w_105_033, w_096_059);
  or2  I165_282(w_165_282, w_053_039, w_090_319);
  nand2 I165_293(w_165_293, w_053_028, w_061_268);
  not1 I165_339(w_165_339, w_066_060);
  or2  I166_021(w_166_021, w_095_038, w_106_176);
  nand2 I166_042(w_166_042, w_034_224, w_107_040);
  and2 I166_075(w_166_075, w_156_115, w_163_187);
  not1 I166_112(w_166_112, w_149_022);
  nand2 I166_181(w_166_181, w_024_027, w_023_024);
  or2  I166_250(w_166_250, w_132_185, w_046_024);
  not1 I166_255(w_166_255, w_161_160);
  or2  I167_011(w_167_011, w_102_030, w_031_061);
  and2 I167_035(w_167_035, w_107_061, w_047_165);
  and2 I167_037(w_167_037, w_032_160, w_131_142);
  nand2 I167_053(w_167_053, w_025_017, w_036_080);
  and2 I167_109(w_167_109, w_105_382, w_053_005);
  not1 I167_136(w_167_136, w_027_178);
  nand2 I167_138(w_167_138, w_049_100, w_056_093);
  nand2 I167_152(w_167_152, w_165_104, w_159_210);
  and2 I167_157(w_167_157, w_122_157, w_018_320);
  and2 I167_168(w_167_168, w_007_062, w_093_276);
  not1 I167_231(w_167_231, w_108_040);
  nand2 I167_302(w_167_302, w_154_013, w_005_211);
  not1 I168_002(w_168_002, w_140_080);
  or2  I168_011(w_168_011, w_127_246, w_120_168);
  or2  I168_015(w_168_015, w_088_421, w_028_255);
  not1 I168_046(w_168_046, w_107_056);
  not1 I168_047(w_168_047, w_076_085);
  not1 I168_053(w_168_053, w_158_000);
  or2  I168_054(w_168_054, w_102_087, w_162_011);
  and2 I168_082(w_168_082, w_029_197, w_162_010);
  not1 I168_103(w_168_103, w_078_136);
  and2 I168_115(w_168_115, w_017_015, w_029_119);
  not1 I168_138(w_168_138, w_086_161);
  nand2 I168_143(w_168_143, w_081_087, w_031_003);
  not1 I168_145(w_168_145, w_157_434);
  not1 I168_151(w_168_151, w_039_241);
  not1 I168_157(w_168_157, w_101_015);
  not1 I169_072(w_169_072, w_083_011);
  or2  I169_215(w_169_215, w_082_197, w_005_173);
  and2 I169_216(w_169_216, w_133_076, w_114_188);
  and2 I169_217(w_169_217, w_141_005, w_024_206);
  and2 I169_222(w_169_222, w_047_164, w_068_036);
  not1 I170_029(w_170_029, w_158_027);
  or2  I170_038(w_170_038, w_015_063, w_032_019);
  not1 I170_061(w_170_061, w_129_000);
  nand2 I170_083(w_170_083, w_049_165, w_022_038);
  or2  I170_089(w_170_089, w_089_138, w_164_058);
  not1 I170_098(w_170_098, w_076_058);
  or2  I170_112(w_170_112, w_075_040, w_110_008);
  not1 I170_137(w_170_137, w_019_041);
  nand2 I170_145(w_170_145, w_120_117, w_096_086);
  nand2 I170_175(w_170_175, w_029_194, w_121_126);
  or2  I170_190(w_170_190, w_162_012, w_149_027);
  nand2 I170_198(w_170_198, w_144_004, w_080_012);
  or2  I170_216(w_170_216, w_025_388, w_021_045);
  nand2 I170_219(w_170_219, w_120_110, w_099_150);
  nand2 I170_221(w_170_221, w_106_354, w_098_010);
  or2  I170_248(w_170_248, w_109_000, w_028_348);
  and2 I171_029(w_171_029, w_078_094, w_085_182);
  and2 I171_084(w_171_084, w_107_032, w_149_011);
  nand2 I171_110(w_171_110, w_006_000, w_037_037);
  nand2 I171_121(w_171_121, w_000_054, w_106_010);
  or2  I171_152(w_171_152, w_034_187, w_096_330);
  and2 I171_173(w_171_173, w_138_215, w_146_061);
  nand2 I171_227(w_171_227, w_089_193, w_051_094);
  nand2 I171_268(w_171_268, w_131_024, w_030_060);
  not1 I171_276(w_171_276, w_103_002);
  not1 I172_009(w_172_009, w_099_111);
  nand2 I172_012(w_172_012, w_063_117, w_171_173);
  and2 I172_018(w_172_018, w_093_115, w_063_206);
  and2 I172_041(w_172_041, w_112_098, w_112_035);
  and2 I172_052(w_172_052, w_068_020, w_136_021);
  nand2 I172_094(w_172_094, w_094_319, w_155_189);
  nand2 I172_102(w_172_102, w_043_063, w_148_129);
  not1 I172_111(w_172_111, w_142_150);
  not1 I172_152(w_172_152, w_066_108);
  not1 I172_168(w_172_168, w_167_035);
  nand2 I172_207(w_172_207, w_045_112, w_093_024);
  and2 I172_224(w_172_224, w_046_056, w_064_003);
  not1 I173_003(w_173_003, w_070_090);
  or2  I173_004(w_173_004, w_129_000, w_026_025);
  or2  I173_062(w_173_062, w_097_163, w_009_094);
  or2  I173_086(w_173_086, w_162_015, w_090_087);
  and2 I173_101(w_173_101, w_145_250, w_033_046);
  nand2 I173_121(w_173_121, w_163_054, w_071_089);
  nand2 I173_134(w_173_134, w_044_307, w_017_098);
  and2 I173_145(w_173_145, w_138_217, w_117_060);
  nand2 I173_204(w_173_204, w_081_053, w_049_060);
  or2  I173_206(w_173_206, w_171_084, w_087_188);
  and2 I173_209(w_173_209, w_042_016, w_153_424);
  nand2 I173_221(w_173_221, w_091_040, w_031_022);
  and2 I173_267(w_173_267, w_127_133, w_008_240);
  nand2 I173_271(w_173_271, w_127_368, w_079_224);
  not1 I173_282(w_173_284, w_173_283);
  not1 I173_283(w_173_285, w_173_284);
  nand2 I173_284(w_173_286, w_064_023, w_173_285);
  or2  I173_285(w_173_287, w_163_330, w_173_286);
  or2  I173_286(w_173_288, w_173_287, w_102_079);
  and2 I173_287(w_173_289, w_007_278, w_173_288);
  and2 I173_288(w_173_290, w_173_289, w_137_021);
  or2  I173_289(w_173_291, w_001_001, w_173_290);
  and2 I173_290(w_173_292, w_173_291, w_046_148);
  and2 I173_291(w_173_283, w_053_006, w_173_292);
  or2  I174_063(w_174_063, w_036_219, w_083_012);
  nand2 I174_090(w_174_090, w_105_116, w_162_014);
  or2  I174_144(w_174_144, w_073_028, w_119_001);
  nand2 I174_147(w_174_147, w_087_004, w_061_190);
  not1 I174_209(w_174_209, w_148_028);
  not1 I174_253(w_174_253, w_080_031);
  not1 I174_278(w_174_278, w_079_407);
  or2  I174_323(w_174_323, w_028_115, w_158_025);
  and2 I174_378(w_174_378, w_124_116, w_008_016);
  or2  I174_399(w_174_399, w_077_123, w_096_018);
  and2 I174_416(w_174_416, w_073_149, w_127_272);
  not1 I174_492(w_174_492, w_009_159);
  nand2 I175_045(w_175_045, w_142_106, w_174_378);
  or2  I175_077(w_175_077, w_069_065, w_002_003);
  nand2 I175_099(w_175_099, w_118_329, w_044_220);
  and2 I175_137(w_175_137, w_086_095, w_115_330);
  and2 I175_171(w_175_171, w_167_136, w_088_012);
  not1 I175_173(w_175_173, w_073_173);
  and2 I175_203(w_175_203, w_028_171, w_073_172);
  nand2 I175_214(w_175_214, w_131_063, w_131_196);
  and2 I175_262(w_175_262, w_065_202, w_074_001);
  nand2 I175_274(w_175_274, w_039_204, w_151_041);
  and2 I175_373(w_175_373, w_152_053, w_015_010);
  not1 I176_036(w_176_036, w_026_104);
  not1 I176_067(w_176_067, w_134_085);
  not1 I176_095(w_176_095, w_014_264);
  not1 I176_111(w_176_111, w_041_036);
  nand2 I176_144(w_176_144, w_032_127, w_071_010);
  or2  I176_196(w_176_196, w_007_092, w_048_020);
  not1 I176_240(w_176_240, w_027_367);
  or2  I176_242(w_176_242, w_134_047, w_074_004);
  nand2 I176_372(w_176_372, w_064_017, w_053_029);
  not1 I176_380(w_176_380, w_012_333);
  and2 I176_383(w_176_383, w_050_015, w_160_025);
  and2 I176_396(w_176_396, w_139_182, w_002_026);
  nand2 I176_397(w_176_397, w_166_112, w_085_055);
  not1 I177_001(w_177_001, w_174_323);
  and2 I177_043(w_177_043, w_119_222, w_155_261);
  not1 I177_089(w_177_089, w_031_051);
  nand2 I177_152(w_177_152, w_155_231, w_084_261);
  and2 I177_212(w_177_212, w_000_000, w_106_003);
  not1 I177_215(w_177_215, w_120_040);
  or2  I177_222(w_177_222, w_018_127, w_147_129);
  or2  I178_029(w_178_029, w_077_125, w_171_121);
  and2 I178_049(w_178_049, w_160_060, w_156_090);
  or2  I178_080(w_178_080, w_019_019, w_067_033);
  and2 I178_104(w_178_104, w_082_113, w_075_109);
  nand2 I178_121(w_178_121, w_073_026, w_003_087);
  not1 I178_172(w_178_172, w_174_399);
  not1 I178_304(w_178_304, w_081_010);
  and2 I178_334(w_178_334, w_061_406, w_149_023);
  or2  I179_002(w_179_002, w_119_101, w_062_005);
  or2  I179_084(w_179_084, w_000_041, w_136_007);
  not1 I179_138(w_179_138, w_123_075);
  or2  I180_007(w_180_007, w_056_056, w_125_081);
  and2 I180_013(w_180_013, w_147_084, w_001_000);
  not1 I180_070(w_180_070, w_128_034);
  not1 I180_120(w_180_120, w_056_026);
  not1 I180_133(w_180_133, w_124_078);
  and2 I180_178(w_180_178, w_103_011, w_057_008);
  nand2 I180_204(w_180_204, w_111_069, w_168_138);
  or2  I180_208(w_180_208, w_012_158, w_031_058);
  or2  I180_210(w_180_210, w_036_163, w_072_054);
  not1 I180_279(w_180_279, w_107_003);
  and2 I181_041(w_181_041, w_108_029, w_116_037);
  or2  I181_047(w_181_047, w_154_058, w_056_169);
  not1 I181_056(w_181_056, w_084_053);
  not1 I181_066(w_181_066, w_079_013);
  or2  I181_073(w_181_073, w_154_106, w_109_001);
  nand2 I181_082(w_181_082, w_062_000, w_109_000);
  not1 I181_087(w_181_087, w_054_074);
  and2 I181_089(w_181_089, w_007_215, w_088_163);
  not1 I181_107(w_181_107, w_154_009);
  and2 I181_119(w_181_119, w_114_080, w_103_002);
  not1 I182_000(w_182_000, w_079_021);
  not1 I182_004(w_182_004, w_006_000);
  or2  I182_010(w_182_010, w_094_003, w_095_058);
  or2  I182_016(w_182_016, w_096_207, w_099_123);
  not1 I182_021(w_182_021, w_044_161);
  and2 I182_024(w_182_024, w_159_158, w_030_199);
  nand2 I182_026(w_182_026, w_047_202, w_112_105);
  nand2 I182_033(w_182_033, w_080_035, w_105_248);
  and2 I182_035(w_182_035, w_008_077, w_028_144);
  nand2 I182_039(w_182_039, w_144_107, w_005_105);
  not1 I182_046(w_182_046, w_031_004);
  and2 I182_059(w_182_059, w_176_372, w_153_186);
  and2 I182_077(w_182_077, w_132_104, w_173_004);
  or2  I182_080(w_182_080, w_034_057, w_123_210);
  and2 I182_087(w_182_087, w_075_094, w_011_093);
  not1 I182_094(w_182_094, w_103_016);
  or2  I182_100(w_182_100, w_014_121, w_033_055);
  and2 I183_019(w_183_019, w_082_002, w_083_177);
  nand2 I183_036(w_183_036, w_164_001, w_051_313);
  or2  I183_038(w_183_038, w_167_168, w_111_028);
  and2 I183_077(w_183_077, w_018_064, w_078_028);
  not1 I184_015(w_184_015, w_091_326);
  and2 I184_021(w_184_021, w_129_000, w_096_010);
  not1 I184_056(w_184_056, w_089_404);
  or2  I184_069(w_184_069, w_009_092, w_153_108);
  and2 I184_095(w_184_095, w_001_000, w_174_416);
  nand2 I184_139(w_184_139, w_010_103, w_008_269);
  and2 I184_158(w_184_158, w_138_122, w_182_004);
  and2 I184_178(w_184_178, w_104_303, w_129_000);
  or2  I184_185(w_184_185, w_143_103, w_121_054);
  nand2 I184_246(w_184_246, w_078_066, w_060_111);
  or2  I184_289(w_184_289, w_180_210, w_030_027);
  and2 I184_368(w_184_368, w_045_210, w_123_062);
  or2  I184_393(w_184_393, w_148_022, w_089_001);
  and2 I184_412(w_184_412, w_113_072, w_023_340);
  or2  I184_418(w_184_418, w_069_012, w_075_122);
  nand2 I184_450(w_184_450, w_025_200, w_119_287);
  not1 I185_031(w_185_031, w_023_256);
  or2  I185_076(w_185_076, w_028_332, w_160_072);
  nand2 I185_109(w_185_109, w_035_069, w_128_015);
  not1 I185_122(w_185_122, w_060_096);
  not1 I185_123(w_185_123, w_164_090);
  not1 I185_126(w_185_126, w_112_150);
  or2  I185_270(w_185_270, w_145_009, w_110_007);
  nand2 I186_008(w_186_008, w_058_073, w_116_116);
  not1 I186_024(w_186_024, w_101_225);
  or2  I186_038(w_186_038, w_076_097, w_065_105);
  nand2 I186_052(w_186_052, w_109_000, w_078_050);
  and2 I186_053(w_186_053, w_092_045, w_014_094);
  or2  I186_056(w_186_056, w_162_013, w_096_024);
  nand2 I186_060(w_186_062, w_186_061, w_080_001);
  and2 I186_061(w_186_063, w_186_062, w_082_144);
  not1 I186_062(w_186_064, w_186_063);
  nand2 I186_063(w_186_065, w_186_064, w_186_085);
  or2  I186_064(w_186_066, w_042_232, w_186_065);
  and2 I186_065(w_186_067, w_052_020, w_186_066);
  not1 I186_066(w_186_068, w_186_067);
  not1 I186_067(w_186_061, w_186_068);
  and2 I186_068(w_186_073, w_186_072, w_093_293);
  nand2 I186_069(w_186_074, w_065_019, w_186_073);
  and2 I186_070(w_186_075, w_001_006, w_186_074);
  or2  I186_071(w_186_076, w_059_211, w_186_075);
  and2 I186_072(w_186_077, w_186_076, w_035_075);
  and2 I186_073(w_186_078, w_186_077, w_108_028);
  or2  I186_074(w_186_079, w_146_011, w_186_078);
  or2  I186_075(w_186_080, w_186_079, w_047_201);
  and2 I186_076(w_186_081, w_162_000, w_186_080);
  and2 I186_077(w_186_082, w_186_081, w_161_219);
  or2  I186_078(w_186_083, w_116_243, w_186_082);
  not1 I186_079(w_186_072, w_186_065);
  and2 I186_080(w_186_085, w_117_279, w_186_083);
  nand2 I187_032(w_187_032, w_071_205, w_080_019);
  not1 I187_053(w_187_053, w_037_121);
  not1 I187_131(w_187_131, w_078_143);
  nand2 I187_155(w_187_155, w_043_141, w_091_077);
  and2 I187_159(w_187_159, w_071_389, w_178_334);
  and2 I188_011(w_188_011, w_033_009, w_007_389);
  not1 I188_034(w_188_034, w_098_023);
  or2  I188_047(w_188_047, w_027_372, w_117_375);
  or2  I188_048(w_188_048, w_140_044, w_155_165);
  nand2 I188_081(w_188_081, w_036_260, w_092_035);
  nand2 I188_089(w_188_089, w_163_007, w_154_075);
  nand2 I188_101(w_188_101, w_025_079, w_122_152);
  or2  I188_105(w_188_105, w_156_153, w_016_374);
  not1 I188_109(w_188_109, w_059_318);
  or2  I189_029(w_189_029, w_166_181, w_153_409);
  and2 I189_058(w_189_058, w_029_096, w_049_065);
  or2  I189_062(w_189_062, w_149_024, w_118_108);
  and2 I189_067(w_189_067, w_025_380, w_147_074);
  and2 I189_135(w_189_135, w_176_067, w_083_105);
  nand2 I189_145(w_189_145, w_048_355, w_080_009);
  and2 I189_213(w_189_213, w_058_051, w_090_079);
  nand2 I189_303(w_189_303, w_177_043, w_137_050);
  or2  I190_014(w_190_014, w_075_099, w_180_279);
  and2 I190_015(w_190_015, w_065_151, w_047_235);
  or2  I190_025(w_190_025, w_028_292, w_085_021);
  and2 I190_027(w_190_027, w_012_340, w_079_453);
  not1 I190_042(w_190_042, w_032_037);
  or2  I190_066(w_190_066, w_122_163, w_151_029);
  or2  I190_077(w_190_077, w_045_115, w_144_062);
  or2  I190_081(w_190_081, w_141_207, w_025_472);
  and2 I190_102(w_190_102, w_130_034, w_134_068);
  nand2 I191_004(w_191_004, w_023_145, w_092_017);
  not1 I191_024(w_191_024, w_067_060);
  and2 I191_075(w_191_075, w_076_097, w_020_072);
  and2 I191_082(w_191_082, w_176_196, w_108_025);
  not1 I191_092(w_191_092, w_088_041);
  and2 I191_150(w_191_150, w_038_054, w_035_005);
  or2  I191_156(w_191_156, w_058_086, w_099_020);
  not1 I191_174(w_191_174, w_123_149);
  not1 I191_181(w_191_181, w_066_067);
  not1 I192_024(w_192_024, w_173_209);
  not1 I192_062(w_192_062, w_082_015);
  and2 I192_086(w_192_086, w_151_033, w_086_068);
  not1 I192_129(w_192_129, w_061_066);
  and2 I192_206(w_192_206, w_033_029, w_025_431);
  not1 I192_221(w_192_221, w_149_018);
  and2 I192_230(w_192_230, w_057_049, w_040_000);
  nand2 I192_247(w_192_247, w_072_097, w_168_082);
  and2 I192_259(w_192_261, w_192_260, w_093_111);
  and2 I192_260(w_192_262, w_192_261, w_187_155);
  and2 I192_261(w_192_263, w_047_173, w_192_262);
  or2  I192_262(w_192_264, w_192_263, w_027_168);
  nand2 I192_263(w_192_265, w_042_212, w_192_264);
  or2  I192_264(w_192_266, w_192_265, w_072_068);
  or2  I192_265(w_192_267, w_192_266, w_142_098);
  nand2 I192_266(w_192_268, w_174_090, w_192_267);
  and2 I192_267(w_192_260, w_192_268, w_117_341);
  and2 I193_012(w_193_012, w_151_036, w_031_037);
  and2 I193_023(w_193_023, w_104_034, w_069_012);
  nand2 I193_039(w_193_039, w_079_304, w_162_010);
  nand2 I193_048(w_193_048, w_180_208, w_043_206);
  or2  I193_082(w_193_082, w_071_156, w_030_133);
  nand2 I194_013(w_194_013, w_053_028, w_109_001);
  and2 I194_058(w_194_058, w_050_173, w_114_146);
  or2  I194_252(w_194_252, w_071_362, w_177_001);
  nand2 I194_259(w_194_259, w_068_011, w_170_219);
  and2 I194_273(w_194_273, w_137_041, w_128_054);
  or2  I195_016(w_195_016, w_014_009, w_061_024);
  not1 I195_041(w_195_041, w_075_070);
  nand2 I195_053(w_195_053, w_159_107, w_024_249);
  nand2 I195_058(w_195_058, w_012_315, w_043_082);
  or2  I195_061(w_195_061, w_080_025, w_118_141);
  not1 I195_076(w_195_076, w_045_090);
  not1 I195_080(w_195_080, w_063_171);
  nand2 I195_081(w_195_081, w_050_067, w_123_124);
  nand2 I195_082(w_195_082, w_128_038, w_092_049);
  nand2 I196_023(w_196_023, w_105_165, w_182_016);
  nand2 I196_069(w_196_069, w_092_068, w_020_098);
  not1 I196_070(w_196_070, w_125_234);
  or2  I196_096(w_196_096, w_148_069, w_142_146);
  nand2 I196_141(w_196_141, w_174_492, w_120_045);
  not1 I196_211(w_196_211, w_192_129);
  and2 I196_214(w_196_214, w_185_076, w_116_137);
  not1 I196_245(w_196_245, w_103_018);
  or2  I196_247(w_196_247, w_175_077, w_142_111);
  and2 I197_024(w_197_024, w_118_046, w_140_266);
  nand2 I197_033(w_197_033, w_123_023, w_151_008);
  or2  I197_081(w_197_081, w_022_053, w_108_045);
  and2 I197_083(w_197_083, w_127_189, w_022_106);
  and2 I197_098(w_197_098, w_058_014, w_078_074);
  not1 I197_102(w_197_102, w_076_013);
  not1 I197_103(w_197_103, w_003_099);
  or2  I197_142(w_197_142, w_143_054, w_050_070);
  nand2 I197_174(w_197_174, w_168_011, w_144_095);
  not1 I197_206(w_197_206, w_052_068);
  or2  I198_020(w_198_020, w_090_163, w_073_222);
  nand2 I198_030(w_198_030, w_109_000, w_038_075);
  and2 I198_071(w_198_071, w_110_060, w_039_270);
  not1 I198_093(w_198_093, w_001_006);
  not1 I198_111(w_198_111, w_176_383);
  and2 I198_179(w_198_179, w_078_067, w_031_046);
  and2 I198_225(w_198_225, w_015_066, w_048_279);
  nand2 I198_323(w_198_323, w_013_163, w_089_273);
  nand2 I198_338(w_198_338, w_195_058, w_150_392);
  nand2 I198_350(w_198_350, w_125_255, w_142_176);
  or2  I199_006(w_199_006, w_123_078, w_077_164);
  and2 I199_007(w_199_007, w_031_053, w_025_258);
  nand2 I199_014(w_199_014, w_076_094, w_051_017);
  nand2 I199_018(w_199_018, w_065_185, w_178_029);
  nand2 I199_019(w_199_019, w_040_004, w_160_132);
  not1 I199_021(w_199_021, w_147_012);
  not1 I199_026(w_199_026, w_161_013);
  not1 I200_011(w_200_011, w_174_209);
  and2 I200_025(w_200_025, w_164_106, w_071_055);
  not1 I200_028(w_200_028, w_137_010);
  nand2 I200_085(w_200_085, w_107_013, w_106_007);
  not1 I200_130(w_200_130, w_136_018);
  and2 I200_186(w_200_186, w_052_104, w_046_004);
  nand2 I200_204(w_200_204, w_086_160, w_126_012);
  nand2 I200_235(w_200_235, w_083_208, w_085_124);
  nand2 I200_253(w_200_253, w_074_001, w_155_237);
  and2 I200_254(w_200_254, w_062_005, w_080_000);
  and2 I201_007(w_201_007, w_098_006, w_063_056);
  not1 I201_017(w_201_017, w_024_064);
  or2  I201_024(w_201_024, w_093_246, w_111_061);
  not1 I201_039(w_201_039, w_088_445);
  and2 I201_090(w_201_090, w_073_191, w_111_005);
  nand2 I201_127(w_201_127, w_047_251, w_178_080);
  not1 I201_196(w_201_196, w_177_215);
  and2 I201_204(w_201_204, w_001_006, w_046_039);
  or2  I201_344(w_201_344, w_066_080, w_093_101);
  nand2 I202_032(w_202_032, w_173_121, w_070_032);
  nand2 I202_056(w_202_056, w_031_013, w_170_145);
  or2  I202_150(w_202_150, w_070_005, w_005_180);
  and2 I202_207(w_202_207, w_005_006, w_039_451);
  not1 I202_230(w_202_230, w_140_026);
  or2  I202_303(w_202_303, w_005_228, w_173_086);
  or2  I202_311(w_202_311, w_119_006, w_088_119);
  or2  I202_411(w_202_411, w_091_052, w_201_204);
  not1 I202_416(w_202_416, w_074_000);
  and2 I203_038(w_203_038, w_176_095, w_190_027);
  not1 I203_055(w_203_055, w_201_017);
  or2  I203_066(w_203_066, w_029_175, w_159_005);
  nand2 I203_071(w_203_071, w_168_015, w_110_095);
  nand2 I203_093(w_203_093, w_193_023, w_022_069);
  nand2 I203_235(w_203_235, w_095_049, w_101_023);
  not1 I203_366(w_203_368, w_203_367);
  or2  I203_367(w_203_369, w_203_390, w_203_368);
  and2 I203_368(w_203_370, w_203_369, w_015_093);
  and2 I203_369(w_203_371, w_203_370, w_035_066);
  and2 I203_370(w_203_372, w_075_103, w_203_371);
  not1 I203_371(w_203_373, w_203_372);
  not1 I203_372(w_203_367, w_203_373);
  not1 I203_373(w_203_378, w_203_377);
  nand2 I203_374(w_203_379, w_203_378, w_005_092);
  and2 I203_375(w_203_380, w_203_379, w_111_081);
  nand2 I203_376(w_203_381, w_203_380, w_015_059);
  and2 I203_377(w_203_382, w_203_381, w_163_054);
  and2 I203_378(w_203_383, w_203_382, w_149_028);
  not1 I203_379(w_203_384, w_203_383);
  not1 I203_380(w_203_385, w_203_384);
  not1 I203_381(w_203_386, w_203_385);
  or2  I203_382(w_203_387, w_203_386, w_011_278);
  nand2 I203_383(w_203_388, w_149_022, w_203_387);
  not1 I203_384(w_203_377, w_203_369);
  and2 I203_385(w_203_390, w_129_000, w_203_388);
  or2  I204_014(w_204_014, w_147_107, w_153_461);
  and2 I204_034(w_204_034, w_033_047, w_195_053);
  or2  I204_058(w_204_058, w_053_011, w_161_031);
  or2  I204_066(w_204_066, w_049_071, w_117_411);
  not1 I204_083(w_204_083, w_019_006);
  not1 I204_117(w_204_117, w_116_208);
  nand2 I204_135(w_204_135, w_072_053, w_170_175);
  not1 I204_223(w_204_223, w_086_055);
  and2 I204_239(w_204_239, w_158_036, w_132_176);
  not1 I204_260(w_204_260, w_189_062);
  and2 I204_274(w_204_274, w_197_103, w_145_219);
  and2 I205_004(w_205_004, w_196_023, w_100_149);
  nand2 I205_007(w_205_007, w_142_000, w_048_265);
  and2 I205_023(w_205_023, w_144_064, w_128_032);
  nand2 I205_047(w_205_047, w_198_179, w_181_082);
  or2  I205_051(w_205_051, w_080_009, w_070_072);
  not1 I205_066(w_205_066, w_001_002);
  not1 I206_030(w_206_030, w_134_075);
  and2 I206_035(w_206_035, w_007_025, w_149_019);
  or2  I206_063(w_206_063, w_070_040, w_006_000);
  and2 I206_098(w_206_098, w_090_089, w_121_269);
  and2 I206_162(w_206_162, w_120_136, w_197_206);
  not1 I206_222(w_206_222, w_029_178);
  nand2 I206_238(w_206_238, w_101_186, w_093_264);
  nand2 I206_331(w_206_331, w_168_011, w_051_246);
  not1 I207_027(w_207_027, w_165_057);
  not1 I207_041(w_207_041, w_182_094);
  nand2 I207_130(w_207_130, w_044_073, w_122_125);
  nand2 I207_204(w_207_204, w_175_045, w_141_061);
  not1 I207_277(w_207_277, w_034_203);
  and2 I207_303(w_207_303, w_100_041, w_172_009);
  nand2 I208_001(w_208_001, w_195_061, w_049_137);
  nand2 I208_004(w_208_004, w_056_131, w_173_003);
  not1 I208_022(w_208_022, w_090_139);
  and2 I208_024(w_208_024, w_127_371, w_104_129);
  not1 I208_032(w_208_032, w_134_069);
  and2 I208_037(w_208_037, w_001_002, w_150_089);
  not1 I208_052(w_208_052, w_153_331);
  and2 I208_076(w_208_076, w_122_110, w_146_050);
  or2  I208_086(w_208_086, w_193_048, w_066_163);
  and2 I208_126(w_208_126, w_070_046, w_122_034);
  not1 I209_033(w_209_033, w_165_028);
  not1 I209_063(w_209_063, w_186_038);
  and2 I209_080(w_209_080, w_019_041, w_049_012);
  or2  I209_129(w_209_129, w_105_041, w_152_022);
  or2  I209_148(w_209_148, w_065_035, w_191_004);
  nand2 I209_406(w_209_406, w_000_083, w_180_204);
  or2  I210_032(w_210_032, w_164_163, w_019_002);
  nand2 I210_060(w_210_060, w_035_040, w_104_002);
  or2  I210_136(w_210_136, w_209_063, w_028_206);
  nand2 I210_140(w_210_140, w_138_013, w_130_142);
  nand2 I210_164(w_210_164, w_127_021, w_170_137);
  nand2 I210_167(w_210_167, w_028_041, w_082_007);
  not1 I210_176(w_210_176, w_191_082);
  not1 I210_212(w_210_212, w_010_451);
  or2  I210_213(w_210_213, w_148_069, w_102_111);
  and2 I210_216(w_210_216, w_102_131, w_144_062);
  nand2 I210_226(w_210_226, w_061_047, w_019_034);
  and2 I210_228(w_210_228, w_110_035, w_004_407);
  or2  I211_055(w_211_055, w_132_133, w_202_056);
  or2  I211_058(w_211_058, w_169_222, w_134_022);
  and2 I211_075(w_211_075, w_196_247, w_176_380);
  and2 I211_077(w_211_077, w_008_058, w_128_031);
  nand2 I211_095(w_211_095, w_069_006, w_019_034);
  or2  I211_118(w_211_118, w_074_000, w_090_228);
  not1 I211_135(w_211_135, w_024_210);
  or2  I211_136(w_211_136, w_140_005, w_200_085);
  not1 I211_257(w_211_257, w_087_039);
  not1 I212_031(w_212_031, w_072_008);
  and2 I212_037(w_212_037, w_067_056, w_210_216);
  or2  I212_052(w_212_052, w_009_086, w_070_090);
  and2 I212_054(w_212_054, w_125_030, w_021_037);
  nand2 I212_063(w_212_063, w_072_020, w_073_133);
  not1 I212_123(w_212_123, w_095_010);
  and2 I212_172(w_212_172, w_171_110, w_101_065);
  and2 I212_192(w_212_192, w_051_023, w_163_035);
  nand2 I213_007(w_213_007, w_096_020, w_103_002);
  or2  I213_014(w_213_014, w_110_156, w_162_009);
  not1 I213_044(w_213_044, w_069_097);
  and2 I213_071(w_213_071, w_148_087, w_000_130);
  not1 I213_177(w_213_177, w_110_020);
  or2  I214_020(w_214_020, w_129_000, w_044_301);
  or2  I214_023(w_214_023, w_001_006, w_153_218);
  and2 I214_026(w_214_026, w_170_061, w_141_163);
  or2  I214_029(w_214_029, w_109_001, w_126_020);
  or2  I214_039(w_214_039, w_166_042, w_181_119);
  nand2 I214_047(w_214_047, w_055_074, w_002_017);
  or2  I214_053(w_214_053, w_068_149, w_148_038);
  nand2 I214_054(w_214_054, w_205_066, w_068_002);
  not1 I214_056(w_214_056, w_204_223);
  not1 I215_008(w_215_008, w_163_210);
  nand2 I215_035(w_215_035, w_159_092, w_063_228);
  not1 I215_054(w_215_054, w_191_092);
  not1 I215_063(w_215_063, w_064_003);
  nand2 I215_075(w_215_075, w_013_050, w_090_128);
  and2 I215_085(w_215_085, w_078_164, w_118_242);
  not1 I215_102(w_215_102, w_058_017);
  nand2 I215_170(w_215_170, w_117_344, w_207_041);
  or2  I215_221(w_215_221, w_066_003, w_032_052);
  nand2 I215_228(w_215_228, w_176_111, w_164_027);
  not1 I215_234(w_215_234, w_041_122);
  and2 I216_003(w_216_003, w_159_128, w_146_161);
  nand2 I216_017(w_216_017, w_050_055, w_158_006);
  and2 I216_041(w_216_041, w_008_241, w_189_303);
  or2  I216_050(w_216_050, w_165_112, w_092_107);
  and2 I216_067(w_216_067, w_068_000, w_083_000);
  and2 I216_072(w_216_072, w_011_196, w_204_135);
  not1 I216_076(w_216_076, w_103_012);
  nand2 I216_123(w_216_123, w_037_132, w_066_126);
  or2  I217_088(w_217_088, w_129_000, w_035_086);
  and2 I217_326(w_217_326, w_060_315, w_202_303);
  nand2 I217_420(w_217_420, w_022_010, w_155_080);
  nand2 I217_423(w_217_423, w_113_041, w_063_028);
  or2  I217_434(w_217_434, w_134_046, w_207_130);
  not1 I218_031(w_218_031, w_195_041);
  not1 I218_048(w_218_048, w_059_018);
  not1 I218_068(w_218_068, w_170_089);
  nand2 I218_081(w_218_081, w_080_004, w_103_013);
  not1 I218_163(w_218_163, w_049_000);
  and2 I218_287(w_218_287, w_180_178, w_140_043);
  not1 I218_396(w_218_396, w_192_024);
  nand2 I219_011(w_219_011, w_060_045, w_092_045);
  or2  I219_041(w_219_041, w_156_225, w_008_064);
  nand2 I219_086(w_219_086, w_109_001, w_168_103);
  and2 I219_220(w_219_220, w_182_021, w_117_362);
  nand2 I219_246(w_219_246, w_060_260, w_196_141);
  or2  I219_254(w_219_254, w_086_100, w_115_423);
  nand2 I219_260(w_219_260, w_190_015, w_101_270);
  nand2 I219_263(w_219_263, w_010_306, w_101_128);
  nand2 I219_290(w_219_290, w_014_038, w_102_149);
  not1 I219_300(w_219_300, w_135_250);
  or2  I219_314(w_219_314, w_067_006, w_086_107);
  and2 I219_361(w_219_361, w_092_023, w_068_149);
  nand2 I220_054(w_220_054, w_136_022, w_031_016);
  nand2 I220_254(w_220_254, w_184_185, w_099_056);
  and2 I220_258(w_220_258, w_098_020, w_213_044);
  nand2 I220_261(w_220_261, w_008_057, w_110_149);
  not1 I220_315(w_220_315, w_010_359);
  nand2 I220_358(w_220_358, w_079_237, w_216_041);
  nand2 I220_440(w_220_440, w_111_014, w_150_225);
  not1 I220_449(w_220_449, w_010_225);
  and2 I220_480(w_220_480, w_097_215, w_150_106);
  and2 I221_012(w_221_012, w_074_005, w_130_021);
  nand2 I221_046(w_221_046, w_184_139, w_111_030);
  or2  I221_050(w_221_050, w_185_270, w_197_174);
  and2 I221_064(w_221_064, w_080_014, w_214_054);
  nand2 I221_079(w_221_079, w_116_023, w_124_031);
  and2 I221_099(w_221_099, w_042_077, w_135_153);
  or2  I221_102(w_221_102, w_058_001, w_101_048);
  and2 I221_107(w_221_107, w_041_013, w_020_009);
  and2 I221_113(w_221_113, w_204_014, w_039_204);
  or2  I222_028(w_222_028, w_043_217, w_210_213);
  and2 I222_030(w_222_030, w_173_271, w_107_068);
  not1 I222_067(w_222_067, w_050_142);
  not1 I222_086(w_222_086, w_085_223);
  not1 I222_100(w_222_100, w_184_289);
  not1 I222_218(w_222_218, w_085_158);
  and2 I222_264(w_222_264, w_030_041, w_026_056);
  not1 I223_066(w_223_066, w_149_004);
  and2 I223_074(w_223_074, w_036_188, w_158_016);
  or2  I223_095(w_223_095, w_016_157, w_182_059);
  nand2 I223_099(w_223_099, w_184_056, w_203_066);
  nand2 I223_168(w_223_168, w_013_007, w_055_037);
  nand2 I223_194(w_223_194, w_075_067, w_090_186);
  or2  I224_000(w_224_000, w_038_058, w_201_039);
  and2 I224_001(w_224_001, w_219_086, w_158_003);
  or2  I224_012(w_224_012, w_000_372, w_028_171);
  or2  I224_016(w_224_016, w_053_014, w_000_314);
  or2  I224_017(w_224_017, w_065_182, w_101_043);
  and2 I224_038(w_224_038, w_022_003, w_215_063);
  not1 I224_045(w_224_045, w_208_024);
  and2 I224_053(w_224_053, w_071_295, w_042_078);
  nand2 I225_005(w_225_005, w_050_175, w_217_326);
  and2 I225_059(w_225_059, w_083_031, w_074_002);
  or2  I225_069(w_225_069, w_114_192, w_216_067);
  or2  I225_167(w_225_167, w_000_381, w_038_026);
  or2  I225_184(w_225_184, w_098_013, w_082_126);
  and2 I225_224(w_225_224, w_196_069, w_210_167);
  or2  I225_248(w_225_248, w_204_034, w_063_024);
  or2  I226_101(w_226_101, w_122_113, w_041_195);
  or2  I226_153(w_226_153, w_206_222, w_018_010);
  and2 I226_188(w_226_188, w_113_052, w_075_080);
  and2 I226_202(w_226_202, w_151_038, w_017_065);
  nand2 I226_310(w_226_310, w_164_012, w_095_094);
  and2 I226_336(w_226_336, w_061_330, w_218_081);
  nand2 I226_395(w_226_397, w_226_396, w_210_060);
  not1 I226_396(w_226_398, w_226_397);
  or2  I226_397(w_226_399, w_040_006, w_226_398);
  not1 I226_398(w_226_400, w_226_399);
  not1 I226_399(w_226_401, w_226_400);
  and2 I226_400(w_226_402, w_226_401, w_200_253);
  and2 I226_401(w_226_403, w_226_402, w_201_007);
  nand2 I226_402(w_226_396, w_226_403, w_169_216);
  or2  I227_019(w_227_019, w_039_343, w_181_066);
  nand2 I227_038(w_227_038, w_215_075, w_026_389);
  nand2 I227_059(w_227_059, w_176_240, w_210_136);
  nand2 I227_061(w_227_061, w_167_231, w_110_149);
  or2  I227_076(w_227_076, w_047_207, w_044_269);
  and2 I227_112(w_227_112, w_058_007, w_172_207);
  not1 I227_150(w_227_150, w_091_254);
  nand2 I227_218(w_227_218, w_095_073, w_186_008);
  nand2 I227_243(w_227_243, w_186_056, w_202_416);
  nand2 I227_285(w_227_285, w_013_017, w_118_175);
  not1 I227_330(w_227_330, w_020_063);
  and2 I228_041(w_228_041, w_103_011, w_094_045);
  not1 I228_066(w_228_066, w_205_007);
  and2 I228_087(w_228_087, w_221_102, w_100_258);
  and2 I228_098(w_228_098, w_106_211, w_052_095);
  not1 I228_284(w_228_284, w_047_422);
  or2  I229_058(w_229_058, w_069_128, w_061_170);
  nand2 I229_092(w_229_092, w_186_053, w_042_077);
  or2  I229_140(w_229_140, w_112_131, w_195_076);
  or2  I229_181(w_229_181, w_162_005, w_102_077);
  or2  I229_269(w_229_269, w_131_191, w_212_054);
  not1 I230_013(w_230_013, w_215_221);
  or2  I230_017(w_230_017, w_124_174, w_207_277);
  nand2 I230_025(w_230_025, w_225_059, w_211_055);
  and2 I230_036(w_230_036, w_214_056, w_184_021);
  nand2 I230_043(w_230_043, w_198_225, w_031_015);
  not1 I230_053(w_230_053, w_068_058);
  nand2 I230_054(w_230_054, w_156_217, w_192_062);
  and2 I231_000(w_231_000, w_028_123, w_017_029);
  and2 I231_005(w_231_005, w_016_339, w_075_056);
  not1 I231_041(w_231_041, w_012_177);
  and2 I231_046(w_231_046, w_099_271, w_184_056);
  and2 I231_049(w_231_049, w_033_042, w_072_065);
  not1 I231_064(w_231_064, w_045_283);
  and2 I231_066(w_231_066, w_038_041, w_220_254);
  nand2 I232_075(w_232_075, w_133_227, w_038_035);
  not1 I233_031(w_233_031, w_217_434);
  and2 I233_065(w_233_065, w_079_065, w_065_093);
  and2 I233_083(w_233_083, w_023_301, w_025_287);
  and2 I233_104(w_233_104, w_227_019, w_034_085);
  and2 I233_203(w_233_203, w_056_177, w_053_027);
  or2  I233_305(w_233_305, w_121_159, w_068_016);
  nand2 I234_001(w_234_001, w_037_068, w_217_420);
  or2  I234_093(w_234_093, w_078_028, w_233_065);
  and2 I234_099(w_234_099, w_019_026, w_013_151);
  not1 I234_115(w_234_115, w_114_153);
  nand2 I234_117(w_234_117, w_048_055, w_172_224);
  nand2 I234_122(w_234_122, w_214_023, w_134_054);
  and2 I235_118(w_235_118, w_075_038, w_107_023);
  or2  I235_211(w_235_211, w_154_078, w_189_135);
  and2 I236_005(w_236_005, w_235_211, w_049_218);
  or2  I236_011(w_236_011, w_016_213, w_093_039);
  not1 I236_018(w_236_018, w_101_019);
  not1 I236_024(w_236_024, w_082_338);
  or2  I236_027(w_236_027, w_212_192, w_225_069);
  nand2 I236_043(w_236_043, w_071_211, w_164_098);
  nand2 I236_046(w_236_046, w_166_250, w_024_111);
  and2 I236_068(w_236_068, w_013_027, w_101_024);
  nand2 I237_008(w_237_008, w_100_163, w_094_010);
  and2 I237_011(w_237_011, w_129_000, w_016_295);
  not1 I237_025(w_237_025, w_003_020);
  not1 I237_037(w_237_037, w_064_044);
  not1 I238_043(w_238_043, w_095_064);
  or2  I238_092(w_238_092, w_182_000, w_042_133);
  nand2 I238_094(w_238_094, w_181_089, w_104_263);
  nand2 I238_126(w_238_126, w_219_254, w_128_043);
  and2 I238_130(w_238_130, w_008_275, w_129_000);
  and2 I238_170(w_238_170, w_233_104, w_189_058);
  and2 I238_190(w_238_190, w_217_088, w_105_426);
  not1 I238_262(w_238_262, w_220_449);
  not1 I238_272(w_238_272, w_122_096);
  not1 I238_309(w_238_309, w_227_285);
  not1 I238_319(w_238_319, w_140_196);
  nand2 I239_017(w_239_017, w_031_001, w_001_001);
  or2  I239_061(w_239_061, w_140_084, w_186_052);
  and2 I239_068(w_239_068, w_023_083, w_021_085);
  not1 I239_092(w_239_092, w_113_035);
  or2  I239_096(w_239_096, w_007_059, w_180_070);
  and2 I239_152(w_239_152, w_114_237, w_236_043);
  not1 I239_236(w_239_236, w_120_140);
  and2 I239_311(w_239_311, w_017_073, w_135_123);
  nand2 I240_026(w_240_026, w_081_038, w_007_230);
  nand2 I240_041(w_240_041, w_148_121, w_083_108);
  nand2 I240_046(w_240_046, w_089_305, w_197_024);
  or2  I240_072(w_240_072, w_184_069, w_062_009);
  or2  I240_122(w_240_122, w_227_330, w_000_490);
  or2  I240_180(w_240_180, w_077_185, w_108_036);
  nand2 I240_182(w_240_182, w_038_089, w_196_245);
  not1 I240_196(w_240_196, w_082_018);
  nand2 I240_206(w_240_206, w_120_136, w_198_350);
  not1 I240_213(w_240_213, w_176_144);
  nand2 I241_014(w_241_014, w_233_083, w_126_016);
  or2  I241_017(w_241_017, w_042_055, w_018_112);
  not1 I241_021(w_241_021, w_219_263);
  and2 I241_047(w_241_047, w_238_130, w_014_093);
  or2  I241_053(w_241_053, w_152_083, w_149_007);
  and2 I241_074(w_241_074, w_123_068, w_071_394);
  or2  I242_038(w_242_038, w_013_120, w_236_046);
  or2  I242_105(w_242_105, w_119_250, w_231_064);
  and2 I242_163(w_242_163, w_216_003, w_093_208);
  not1 I242_346(w_242_346, w_004_274);
  nand2 I243_190(w_243_190, w_061_130, w_005_192);
  not1 I244_022(w_244_022, w_086_149);
  and2 I244_075(w_244_075, w_223_074, w_240_046);
  or2  I244_089(w_244_089, w_052_097, w_145_393);
  or2  I244_109(w_244_109, w_169_072, w_188_081);
  or2  I244_135(w_244_135, w_228_098, w_201_090);
  not1 I244_160(w_244_160, w_116_029);
  not1 I245_019(w_245_019, w_016_212);
  not1 I245_057(w_245_057, w_030_012);
  not1 I245_106(w_245_106, w_036_067);
  not1 I245_118(w_245_118, w_152_147);
  or2  I245_121(w_245_121, w_011_057, w_111_087);
  nand2 I245_135(w_245_135, w_170_248, w_142_086);
  not1 I245_193(w_245_193, w_022_149);
  not1 I246_019(w_246_019, w_165_092);
  not1 I246_065(w_246_065, w_166_255);
  or2  I246_078(w_246_078, w_226_188, w_060_344);
  and2 I246_093(w_246_093, w_101_126, w_149_026);
  not1 I246_258(w_246_258, w_200_025);
  not1 I246_273(w_246_273, w_134_043);
  and2 I246_363(w_246_363, w_177_152, w_088_031);
  nand2 I247_040(w_247_040, w_004_014, w_116_028);
  or2  I247_054(w_247_054, w_025_174, w_050_051);
  and2 I247_065(w_247_065, w_215_008, w_168_143);
  nand2 I247_223(w_247_223, w_171_152, w_114_040);
  not1 I247_230(w_247_230, w_130_072);
  nand2 I247_254(w_247_254, w_075_121, w_060_040);
  and2 I248_029(w_248_029, w_155_101, w_040_005);
  and2 I248_115(w_248_115, w_007_244, w_229_269);
  nand2 I248_133(w_248_133, w_238_319, w_243_190);
  or2  I248_243(w_248_243, w_053_006, w_117_201);
  nand2 I248_360(w_248_360, w_053_034, w_239_096);
  and2 I249_029(w_249_029, w_144_010, w_238_309);
  not1 I249_031(w_249_031, w_246_258);
  or2  I249_033(w_249_033, w_159_055, w_247_054);
  not1 I249_052(w_249_052, w_125_117);
  and2 I249_068(w_249_068, w_011_012, w_033_014);
  or2  I249_082(w_249_082, w_098_014, w_220_258);
  or2  I249_083(w_249_083, w_108_032, w_034_016);
  and2 I249_089(w_249_089, w_185_109, w_093_318);
  and2 I249_102(w_249_102, w_215_170, w_020_052);
  or2  I250_002(w_250_002, w_153_007, w_211_058);
  not1 I250_029(w_250_029, w_136_017);
  nand2 I250_035(w_250_035, w_182_026, w_050_113);
  or2  I250_044(w_250_044, w_031_018, w_117_410);
  or2  I250_047(w_250_047, w_073_176, w_210_140);
  not1 I250_049(w_250_049, w_021_051);
  or2  I250_057(w_250_057, w_055_039, w_239_311);
  not1 I251_017(w_251_017, w_017_141);
  nand2 I251_038(w_251_038, w_034_014, w_184_450);
  nand2 I251_056(w_251_056, w_146_017, w_019_027);
  and2 I251_085(w_251_085, w_084_010, w_046_004);
  not1 I251_098(w_251_098, w_227_218);
  not1 I251_112(w_251_112, w_249_089);
  not1 I251_113(w_251_113, w_201_344);
  or2  I251_124(w_251_124, w_103_012, w_017_064);
  not1 I252_002(w_252_002, w_227_059);
  nand2 I252_041(w_252_041, w_025_023, w_062_003);
  or2  I252_092(w_252_092, w_184_158, w_107_043);
  and2 I252_147(w_252_147, w_157_393, w_017_136);
  and2 I252_234(w_252_234, w_122_128, w_012_119);
  or2  I252_279(w_252_279, w_091_326, w_183_019);
  and2 I252_327(w_252_327, w_027_041, w_146_041);
  and2 I252_383(w_252_383, w_152_191, w_142_083);
  and2 I253_010(w_253_010, w_103_005, w_160_013);
  nand2 I253_023(w_253_023, w_246_019, w_153_255);
  nand2 I253_048(w_253_048, w_014_226, w_171_029);
  and2 I253_097(w_253_097, w_190_042, w_173_101);
  or2  I253_123(w_253_123, w_032_074, w_199_018);
  nand2 I253_140(w_253_140, w_010_063, w_041_037);
  not1 I254_014(w_254_014, w_140_110);
  not1 I254_037(w_254_037, w_046_035);
  nand2 I254_050(w_254_050, w_003_061, w_246_093);
  and2 I254_101(w_254_101, w_034_097, w_185_126);
  or2  I255_037(w_255_037, w_132_113, w_131_041);
  nand2 I255_057(w_255_057, w_099_277, w_253_123);
  nand2 I255_068(w_255_068, w_039_356, w_084_055);
  and2 I255_186(w_255_186, w_061_117, w_157_019);
  not1 I255_197(w_255_197, w_024_165);
  or2  I256_005(w_256_005, w_154_103, w_120_016);
  or2  I256_011(w_256_011, w_145_073, w_083_171);
  and2 I256_072(w_256_072, w_164_119, w_161_141);
  not1 I256_125(w_256_125, w_106_359);
  nand2 I256_134(w_256_134, w_106_168, w_180_007);
  not1 I257_014(w_257_014, w_092_038);
  and2 I257_040(w_257_040, w_063_139, w_102_127);
  not1 I257_048(w_257_048, w_049_403);
  or2  I257_050(w_257_050, w_184_412, w_255_186);
  and2 I257_052(w_257_052, w_145_009, w_106_202);
  nand2 I257_073(w_257_073, w_116_275, w_145_063);
  or2  I257_102(w_257_102, w_254_014, w_118_054);
  and2 I257_168(w_257_168, w_037_047, w_191_156);
  not1 I257_213(w_257_213, w_003_075);
  nand2 I257_214(w_257_214, w_193_012, w_059_223);
  nand2 I258_022(w_258_022, w_047_013, w_039_494);
  and2 I258_045(w_258_045, w_099_013, w_184_246);
  nand2 I258_046(w_258_046, w_017_061, w_097_182);
  or2  I258_190(w_258_190, w_214_020, w_056_149);
  and2 I258_261(w_258_261, w_081_004, w_222_086);
  and2 I259_042(w_259_042, w_247_040, w_250_057);
  not1 I259_044(w_259_044, w_058_038);
  not1 I259_079(w_259_079, w_150_176);
  not1 I259_102(w_259_102, w_204_058);
  nand2 I259_104(w_259_104, w_134_042, w_159_007);
  or2  I259_131(w_259_131, w_054_134, w_110_094);
  or2  I259_153(w_259_153, w_055_064, w_035_071);
  or2  I260_000(w_260_000, w_034_202, w_131_141);
  and2 I260_054(w_260_054, w_133_232, w_092_073);
  or2  I260_057(w_260_057, w_047_322, w_214_023);
  not1 I260_063(w_260_063, w_103_004);
  or2  I260_074(w_260_074, w_210_164, w_155_110);
  not1 I260_076(w_260_076, w_184_095);
  nand2 I260_163(w_260_163, w_104_112, w_011_268);
  nand2 I260_181(w_260_181, w_122_092, w_024_139);
  or2  I261_041(w_261_041, w_162_008, w_188_101);
  not1 I261_083(w_261_083, w_155_072);
  or2  I261_115(w_261_115, w_166_075, w_027_201);
  nand2 I262_050(w_262_050, w_251_038, w_209_129);
  or2  I262_062(w_262_064, w_262_063, w_073_036);
  or2  I262_063(w_262_065, w_250_002, w_262_064);
  or2  I262_064(w_262_066, w_211_257, w_262_065);
  and2 I262_065(w_262_067, w_106_395, w_262_066);
  or2  I262_066(w_262_068, w_262_067, w_164_136);
  not1 I262_067(w_262_069, w_262_068);
  or2  I262_068(w_262_070, w_262_069, w_129_000);
  and2 I262_069(w_262_071, w_252_327, w_262_070);
  not1 I262_070(w_262_072, w_262_071);
  and2 I262_071(w_262_073, w_262_072, w_250_047);
  and2 I262_072(w_262_074, w_139_176, w_262_073);
  and2 I262_073(w_262_063, w_121_034, w_262_074);
  nand2 I263_020(w_263_020, w_072_086, w_015_031);
  nand2 I263_026(w_263_026, w_219_314, w_072_045);
  and2 I263_040(w_263_040, w_032_187, w_222_264);
  not1 I263_053(w_263_053, w_133_282);
  not1 I263_114(w_263_114, w_198_030);
  not1 I263_194(w_263_194, w_033_004);
  and2 I264_012(w_264_012, w_089_101, w_120_061);
  or2  I264_064(w_264_064, w_113_039, w_153_025);
  not1 I264_085(w_264_085, w_212_063);
  nand2 I264_125(w_264_125, w_122_141, w_219_041);
  not1 I264_191(w_264_191, w_150_334);
  or2  I264_275(w_264_275, w_067_050, w_047_001);
  not1 I264_355(w_264_355, w_200_011);
  and2 I265_000(w_265_000, w_124_147, w_112_074);
  and2 I265_003(w_265_003, w_214_047, w_108_046);
  nand2 I265_006(w_265_006, w_252_002, w_113_030);
  not1 I265_017(w_265_017, w_200_254);
  nand2 I266_076(w_266_076, w_095_017, w_063_076);
  nand2 I266_111(w_266_111, w_233_305, w_106_271);
  nand2 I266_314(w_266_314, w_162_011, w_100_193);
  or2  I266_408(w_266_408, w_108_000, w_198_020);
  nand2 I267_128(w_267_128, w_152_134, w_024_230);
  nand2 I267_222(w_267_222, w_199_014, w_244_075);
  not1 I267_355(w_267_355, w_227_243);
  and2 I267_389(w_267_389, w_103_003, w_228_041);
  not1 I268_018(w_268_018, w_036_094);
  or2  I268_025(w_268_025, w_162_001, w_002_021);
  not1 I268_040(w_268_040, w_120_110);
  or2  I268_139(w_268_139, w_202_311, w_094_062);
  or2  I268_150(w_268_150, w_103_017, w_172_009);
  and2 I269_029(w_269_029, w_152_132, w_162_014);
  and2 I269_038(w_269_038, w_160_138, w_048_347);
  and2 I269_043(w_269_043, w_055_046, w_146_037);
  or2  I269_055(w_269_055, w_157_165, w_205_004);
  not1 I269_059(w_269_059, w_045_009);
  or2  I270_021(w_270_021, w_198_071, w_167_109);
  or2  I270_054(w_270_054, w_051_104, w_151_007);
  nand2 I270_111(w_270_111, w_168_145, w_121_242);
  nand2 I270_190(w_270_190, w_018_259, w_015_073);
  and2 I270_255(w_270_255, w_069_008, w_108_050);
  nand2 I271_026(w_271_026, w_088_315, w_151_038);
  and2 I271_048(w_271_048, w_038_044, w_102_031);
  and2 I271_118(w_271_118, w_085_244, w_083_103);
  and2 I271_151(w_271_151, w_160_114, w_259_044);
  not1 I271_172(w_271_172, w_103_000);
  or2  I271_254(w_271_254, w_201_024, w_122_045);
  not1 I271_280(w_271_280, w_153_125);
  and2 I271_338(w_271_338, w_149_000, w_199_018);
  nand2 I272_003(w_272_003, w_057_028, w_208_086);
  not1 I272_009(w_272_009, w_170_221);
  or2  I272_010(w_272_010, w_099_223, w_093_072);
  and2 I272_019(w_272_019, w_093_110, w_152_059);
  and2 I272_020(w_272_020, w_211_077, w_251_112);
  nand2 I272_022(w_272_022, w_182_033, w_119_282);
  nand2 I272_024(w_272_024, w_005_023, w_123_026);
  nand2 I272_029(w_272_029, w_200_204, w_175_173);
  or2  I272_031(w_272_031, w_119_157, w_089_307);
  not1 I273_023(w_273_023, w_188_034);
  nand2 I273_044(w_273_044, w_152_029, w_135_113);
  or2  I273_071(w_273_071, w_049_388, w_073_111);
  and2 I273_142(w_273_142, w_003_032, w_143_099);
  or2  I273_143(w_273_143, w_110_193, w_117_322);
  not1 I274_017(w_274_017, w_064_018);
  not1 I274_034(w_274_034, w_265_000);
  nand2 I274_149(w_274_149, w_195_058, w_103_012);
  and2 I274_192(w_274_192, w_134_034, w_257_213);
  not1 I275_053(w_275_053, w_257_102);
  and2 I275_054(w_275_054, w_069_149, w_046_060);
  or2  I275_088(w_275_088, w_104_014, w_218_048);
  or2  I275_097(w_275_097, w_132_067, w_028_129);
  nand2 I275_117(w_275_117, w_081_088, w_052_007);
  and2 I275_123(w_275_123, w_123_188, w_044_154);
  and2 I276_117(w_276_117, w_045_284, w_024_205);
  nand2 I277_003(w_277_003, w_179_002, w_082_275);
  and2 I277_005(w_277_005, w_061_027, w_028_381);
  or2  I277_013(w_277_013, w_258_045, w_016_136);
  not1 I277_015(w_277_015, w_095_091);
  not1 I277_046(w_277_046, w_006_000);
  or2  I278_079(w_278_079, w_028_356, w_117_261);
  or2  I278_118(w_278_118, w_010_170, w_148_251);
  nand2 I279_071(w_279_071, w_095_014, w_253_097);
  or2  I279_309(w_279_309, w_177_089, w_008_148);
  or2  I279_345(w_279_345, w_197_033, w_005_252);
  not1 I279_415(w_279_415, w_134_026);
  or2  I280_008(w_280_008, w_210_228, w_227_038);
  or2  I280_025(w_280_025, w_115_171, w_125_186);
  or2  I280_060(w_280_060, w_011_072, w_117_238);
  and2 I280_063(w_280_063, w_249_082, w_226_153);
  and2 I281_002(w_281_002, w_100_301, w_011_130);
  or2  I281_009(w_281_009, w_128_031, w_154_047);
  nand2 I281_010(w_281_010, w_067_032, w_065_036);
  nand2 I281_015(w_281_015, w_143_092, w_259_104);
  and2 I281_016(w_281_016, w_162_017, w_081_069);
  not1 I282_037(w_282_037, w_220_440);
  not1 I282_046(w_282_046, w_135_203);
  not1 I282_065(w_282_065, w_024_081);
  nand2 I282_096(w_282_096, w_004_425, w_275_097);
  and2 I282_122(w_282_122, w_241_074, w_055_079);
  and2 I283_026(w_283_026, w_077_029, w_143_002);
  and2 I283_139(w_283_139, w_244_160, w_047_367);
  and2 I283_169(w_283_169, w_100_402, w_001_004);
  or2  I283_188(w_283_188, w_115_424, w_203_071);
  not1 I283_224(w_283_224, w_080_012);
  or2  I284_013(w_284_013, w_239_061, w_004_442);
  or2  I284_122(w_284_122, w_173_204, w_267_355);
  and2 I284_265(w_284_265, w_156_066, w_027_339);
  or2  I285_000(w_285_000, w_120_009, w_000_040);
  or2  I285_018(w_285_018, w_228_087, w_182_035);
  or2  I285_021(w_285_021, w_169_215, w_277_013);
  and2 I285_022(w_285_022, w_206_238, w_013_200);
  not1 I285_024(w_285_026, w_285_025);
  not1 I285_025(w_285_027, w_285_026);
  nand2 I285_026(w_285_028, w_285_027, w_042_206);
  or2  I285_027(w_285_029, w_285_028, w_197_081);
  and2 I285_028(w_285_030, w_087_281, w_285_029);
  nand2 I285_029(w_285_031, w_285_030, w_260_181);
  and2 I285_030(w_285_032, w_285_031, w_045_276);
  or2  I285_031(w_285_033, w_178_304, w_285_032);
  or2  I285_032(w_285_034, w_129_000, w_285_033);
  or2  I285_033(w_285_035, w_285_034, w_017_071);
  or2  I285_034(w_285_025, w_098_011, w_285_035);
  or2  I286_002(w_286_002, w_010_162, w_221_012);
  nand2 I286_039(w_286_039, w_129_000, w_189_145);
  and2 I286_054(w_286_054, w_245_118, w_078_062);
  and2 I286_088(w_286_088, w_039_254, w_265_017);
  and2 I286_234(w_286_234, w_163_383, w_079_040);
  or2  I286_434(w_286_434, w_097_164, w_032_124);
  not1 I287_000(w_287_000, w_285_021);
  nand2 I287_135(w_287_135, w_211_095, w_065_219);
  not1 I287_179(w_287_179, w_054_088);
  or2  I287_254(w_287_254, w_216_050, w_034_196);
  nand2 I287_256(w_287_256, w_244_022, w_108_043);
  or2  I287_308(w_287_308, w_181_087, w_283_188);
  and2 I287_423(w_287_423, w_264_355, w_014_018);
  and2 I287_477(w_287_477, w_052_038, w_108_056);
  nand2 I288_027(w_288_027, w_199_026, w_122_002);
  and2 I288_190(w_288_190, w_048_247, w_222_100);
  or2  I289_079(w_289_079, w_267_128, w_150_320);
  or2  I289_089(w_289_089, w_249_068, w_021_076);
  not1 I289_097(w_289_097, w_047_030);
  not1 I289_099(w_289_099, w_254_050);
  nand2 I289_118(w_289_118, w_136_007, w_136_029);
  or2  I289_120(w_289_120, w_095_017, w_236_027);
  not1 I289_124(w_289_124, w_054_084);
  and2 I290_019(w_290_019, w_251_098, w_021_002);
  nand2 I290_069(w_290_069, w_111_088, w_048_061);
  not1 I291_015(w_291_015, w_136_019);
  and2 I291_122(w_291_122, w_238_094, w_268_150);
  not1 I291_131(w_291_131, w_083_098);
  and2 I292_087(w_292_087, w_061_041, w_218_068);
  not1 I292_099(w_292_099, w_280_060);
  or2  I292_106(w_292_106, w_111_061, w_266_111);
  nand2 I293_011(w_293_011, w_216_076, w_240_196);
  nand2 I293_037(w_293_037, w_286_234, w_128_013);
  not1 I293_099(w_293_099, w_096_004);
  and2 I293_134(w_293_134, w_176_242, w_258_261);
  nand2 I294_001(w_294_001, w_151_010, w_204_083);
  or2  I294_037(w_294_037, w_134_002, w_030_116);
  and2 I294_111(w_294_111, w_060_370, w_114_102);
  not1 I294_185(w_294_185, w_034_166);
  and2 I295_050(w_295_050, w_058_074, w_241_053);
  not1 I295_090(w_295_090, w_079_320);
  nand2 I295_171(w_295_171, w_237_037, w_091_354);
  or2  I295_208(w_295_208, w_154_050, w_012_324);
  not1 I295_315(w_295_315, w_093_064);
  nand2 I296_135(w_296_135, w_238_092, w_152_062);
  nand2 I296_144(w_296_144, w_069_108, w_231_046);
  and2 I296_401(w_296_401, w_146_087, w_281_002);
  nand2 I296_411(w_296_411, w_252_041, w_034_129);
  not1 I297_016(w_297_016, w_003_027);
  not1 I297_021(w_297_021, w_191_174);
  not1 I297_027(w_297_027, w_030_184);
  or2  I297_038(w_297_038, w_163_156, w_020_023);
  nand2 I297_287(w_297_287, w_263_114, w_040_002);
  not1 I297_365(w_297_365, w_092_009);
  nand2 I298_024(w_298_024, w_151_023, w_271_026);
  or2  I298_031(w_298_031, w_264_275, w_245_057);
  and2 I298_112(w_298_112, w_139_016, w_255_197);
  or2  I298_179(w_298_179, w_056_162, w_121_247);
  and2 I298_191(w_298_191, w_224_016, w_218_287);
  nand2 I299_032(w_299_032, w_155_322, w_209_406);
  and2 I300_121(w_300_121, w_052_034, w_275_117);
  not1 I300_202(w_300_202, w_287_254);
  not1 I300_233(w_300_233, w_212_172);
  nand2 I300_250(w_300_250, w_201_127, w_147_106);
  or2  I301_027(w_301_027, w_143_018, w_253_010);
  nand2 I301_161(w_301_161, w_017_047, w_241_014);
  and2 I302_029(w_302_029, w_042_044, w_240_182);
  and2 I302_079(w_302_079, w_033_047, w_022_110);
  not1 I302_097(w_302_097, w_198_111);
  or2  I302_103(w_302_103, w_297_287, w_084_086);
  nand2 I303_011(w_303_011, w_269_029, w_241_047);
  nand2 I303_084(w_303_084, w_026_189, w_074_003);
  not1 I303_127(w_303_127, w_272_019);
  not1 I303_144(w_303_144, w_009_004);
  not1 I303_162(w_303_162, w_252_234);
  or2  I303_178(w_303_178, w_302_079, w_027_009);
  nand2 I303_196(w_303_198, w_303_215, w_303_197);
  not1 I303_197(w_303_199, w_303_198);
  and2 I303_198(w_303_200, w_153_093, w_303_199);
  not1 I303_199(w_303_197, w_303_200);
  not1 I303_200(w_303_205, w_303_204);
  not1 I303_201(w_303_206, w_303_205);
  or2  I303_202(w_303_207, w_303_206, w_115_346);
  nand2 I303_203(w_303_208, w_303_207, w_239_017);
  not1 I303_204(w_303_209, w_303_208);
  and2 I303_205(w_303_210, w_303_209, w_277_046);
  not1 I303_206(w_303_211, w_303_210);
  and2 I303_207(w_303_212, w_181_107, w_303_211);
  or2  I303_208(w_303_213, w_303_212, w_106_146);
  not1 I303_209(w_303_204, w_303_198);
  and2 I303_210(w_303_215, w_040_004, w_303_213);
  and2 I304_065(w_304_065, w_213_007, w_289_079);
  or2  I304_136(w_304_136, w_112_028, w_265_006);
  not1 I304_188(w_304_188, w_223_066);
  or2  I305_007(w_305_007, w_211_136, w_270_021);
  nand2 I305_054(w_305_054, w_198_338, w_285_000);
  and2 I305_057(w_305_057, w_176_036, w_172_111);
  and2 I305_085(w_305_085, w_061_376, w_209_080);
  nand2 I306_004(w_306_004, w_149_005, w_289_099);
  and2 I306_007(w_306_007, w_217_423, w_042_111);
  not1 I306_088(w_306_088, w_231_005);
  not1 I306_287(w_306_287, w_023_177);
  nand2 I307_002(w_307_002, w_122_026, w_122_114);
  and2 I307_062(w_307_062, w_116_108, w_125_166);
  and2 I307_075(w_307_075, w_015_022, w_142_070);
  nand2 I307_123(w_307_123, w_239_152, w_182_080);
  or2  I307_129(w_307_129, w_032_052, w_157_229);
  nand2 I307_183(w_307_183, w_141_154, w_266_408);
  nand2 I308_024(w_308_024, w_035_100, w_011_127);
  or2  I308_027(w_308_027, w_133_357, w_059_478);
  or2  I308_050(w_308_050, w_020_156, w_156_302);
  or2  I309_026(w_309_026, w_143_070, w_281_009);
  not1 I309_065(w_309_065, w_262_050);
  nand2 I309_073(w_309_073, w_154_062, w_297_365);
  and2 I309_095(w_309_095, w_284_013, w_074_004);
  and2 I309_115(w_309_115, w_094_416, w_036_209);
  or2  I309_145(w_309_145, w_261_041, w_031_051);
  nand2 I310_070(w_310_070, w_114_015, w_085_159);
  nand2 I310_071(w_310_071, w_098_018, w_192_247);
  and2 I310_072(w_310_072, w_196_214, w_073_181);
  or2  I310_184(w_310_184, w_056_076, w_257_073);
  nand2 I310_226(w_310_226, w_221_107, w_185_123);
  or2  I311_067(w_311_067, w_112_078, w_222_028);
  nand2 I311_134(w_311_134, w_282_046, w_119_141);
  or2  I311_149(w_311_149, w_199_021, w_225_167);
  nand2 I311_174(w_311_174, w_187_159, w_104_385);
  nand2 I312_068(w_312_068, w_300_233, w_192_230);
  and2 I312_123(w_312_123, w_004_247, w_247_223);
  not1 I312_137(w_312_137, w_026_017);
  not1 I312_171(w_312_171, w_068_099);
  and2 I312_174(w_312_174, w_103_005, w_295_050);
  nand2 I312_199(w_312_199, w_223_168, w_095_084);
  or2  I312_222(w_312_222, w_139_025, w_061_025);
  nand2 I313_074(w_313_074, w_117_406, w_306_007);
  nand2 I313_089(w_313_089, w_197_102, w_063_113);
  and2 I313_092(w_313_092, w_275_123, w_208_032);
  nand2 I313_111(w_313_111, w_012_322, w_182_039);
  nand2 I313_119(w_313_119, w_233_031, w_277_003);
  nand2 I313_151(w_313_151, w_220_480, w_003_062);
  nand2 I314_093(w_314_093, w_309_026, w_096_127);
  not1 I314_142(w_314_142, w_151_021);
  and2 I314_214(w_314_214, w_106_286, w_092_014);
  and2 I314_369(w_314_369, w_180_120, w_312_068);
  or2  I314_382(w_314_382, w_093_000, w_155_329);
  not1 I315_122(w_315_122, w_067_004);
  nand2 I315_242(w_315_242, w_205_051, w_063_022);
  not1 I315_288(w_315_288, w_236_011);
  not1 I315_325(w_315_325, w_113_045);
  or2  I316_014(w_316_014, w_074_004, w_101_074);
  and2 I316_021(w_316_021, w_126_005, w_266_076);
  or2  I316_044(w_316_044, w_137_054, w_264_012);
  nand2 I316_046(w_316_046, w_002_025, w_225_224);
  and2 I316_057(w_316_057, w_210_212, w_002_006);
  or2  I316_224(w_316_224, w_073_218, w_024_106);
  and2 I317_116(w_317_116, w_182_046, w_130_037);
  or2  I317_248(w_317_248, w_006_000, w_068_129);
  and2 I317_304(w_317_304, w_103_007, w_101_301);
  and2 I317_340(w_317_342, w_119_107, w_317_341);
  not1 I317_341(w_317_343, w_317_342);
  or2  I317_342(w_317_344, w_317_343, w_313_092);
  or2  I317_343(w_317_345, w_317_344, w_234_117);
  nand2 I317_344(w_317_346, w_225_184, w_317_345);
  nand2 I317_345(w_317_347, w_298_179, w_317_346);
  nand2 I317_346(w_317_348, w_317_347, w_109_001);
  not1 I317_347(w_317_349, w_317_348);
  or2  I317_348(w_317_350, w_099_267, w_317_349);
  or2  I317_349(w_317_351, w_317_350, w_206_098);
  and2 I317_350(w_317_341, w_317_351, w_079_170);
  or2  I318_049(w_318_049, w_246_065, w_215_085);
  and2 I318_084(w_318_084, w_259_079, w_036_152);
  and2 I318_159(w_318_159, w_130_012, w_116_038);
  and2 I318_290(w_318_290, w_227_076, w_108_050);
  and2 I318_309(w_318_309, w_113_056, w_184_368);
  not1 I318_342(w_318_342, w_308_050);
  not1 I318_382(w_318_383, w_318_382);
  not1 I318_383(w_318_384, w_318_383);
  and2 I318_384(w_318_385, w_318_384, w_318_401);
  or2  I318_385(w_318_386, w_066_014, w_318_385);
  and2 I318_386(w_318_387, w_318_386, w_173_145);
  and2 I318_387(w_318_388, w_318_387, w_213_014);
  not1 I318_388(w_318_389, w_318_388);
  or2  I318_389(w_318_390, w_180_013, w_318_389);
  not1 I318_390(w_318_382, w_318_390);
  or2  I318_391(w_318_395, w_178_172, w_318_394);
  not1 I318_392(w_318_396, w_318_395);
  and2 I318_393(w_318_397, w_318_396, w_147_151);
  nand2 I318_394(w_318_398, w_020_085, w_318_397);
  or2  I318_395(w_318_399, w_318_398, w_023_264);
  not1 I318_396(w_318_394, w_318_385);
  and2 I318_397(w_318_401, w_135_049, w_318_399);
  and2 I319_007(w_319_007, w_007_272, w_170_216);
  or2  I319_030(w_319_030, w_125_463, w_052_018);
  not1 I319_064(w_319_064, w_016_070);
  nand2 I319_081(w_319_081, w_064_035, w_163_016);
  nand2 I319_099(w_319_099, w_230_036, w_233_203);
  nand2 I320_108(w_320_108, w_005_157, w_237_008);
  or2  I320_219(w_320_219, w_050_043, w_312_123);
  not1 I320_260(w_320_260, w_297_021);
  nand2 I321_001(w_321_001, w_117_138, w_161_261);
  and2 I321_056(w_321_056, w_237_011, w_216_072);
  or2  I321_096(w_321_096, w_108_050, w_151_000);
  or2  I321_108(w_321_108, w_302_097, w_247_065);
  and2 I322_007(w_322_007, w_199_007, w_024_055);
  not1 I322_030(w_322_030, w_197_098);
  nand2 I323_000(w_323_000, w_017_051, w_018_111);
  nand2 I323_003(w_323_003, w_172_152, w_020_165);
  not1 I323_033(w_323_033, w_319_007);
  and2 I323_046(w_323_046, w_203_093, w_022_037);
  not1 I323_057(w_323_057, w_172_102);
  nand2 I324_047(w_324_047, w_115_314, w_093_258);
  or2  I325_126(w_325_126, w_152_056, w_067_062);
  not1 I325_190(w_325_190, w_039_093);
  and2 I325_206(w_325_206, w_040_004, w_125_249);
  and2 I325_464(w_325_464, w_074_002, w_252_383);
  nand2 I326_028(w_326_028, w_323_003, w_220_315);
  not1 I326_035(w_326_035, w_047_137);
  not1 I326_040(w_326_040, w_245_135);
  and2 I326_053(w_326_053, w_038_021, w_264_191);
  not1 I326_069(w_326_069, w_073_017);
  nand2 I327_041(w_327_041, w_044_151, w_093_053);
  and2 I327_163(w_327_163, w_041_208, w_117_403);
  or2  I327_172(w_327_172, w_181_041, w_281_015);
  or2  I327_176(w_327_176, w_004_402, w_009_038);
  and2 I328_038(w_328_038, w_327_172, w_100_219);
  or2  I328_058(w_328_058, w_040_000, w_280_025);
  nand2 I328_215(w_328_215, w_120_109, w_200_028);
  and2 I328_241(w_328_241, w_184_418, w_302_103);
  not1 I328_297(w_328_297, w_094_229);
  not1 I328_459(w_328_459, w_182_010);
  nand2 I329_074(w_329_074, w_273_023, w_068_103);
  or2  I329_237(w_329_237, w_260_054, w_152_120);
  or2  I329_287(w_329_287, w_025_322, w_112_020);
  not1 I329_321(w_329_321, w_125_359);
  not1 I329_342(w_329_342, w_069_040);
  not1 I329_431(w_329_431, w_300_202);
  nand2 I330_029(w_330_029, w_190_102, w_087_061);
  not1 I330_134(w_330_134, w_022_025);
  and2 I330_154(w_330_154, w_295_315, w_176_397);
  and2 I330_364(w_330_364, w_251_085, w_004_105);
  and2 I331_017(w_331_017, w_215_035, w_249_083);
  or2  I331_022(w_331_022, w_175_137, w_191_181);
  not1 I331_032(w_331_032, w_252_147);
  and2 I331_042(w_331_042, w_067_008, w_130_171);
  and2 I332_014(w_332_014, w_100_215, w_014_188);
  or2  I332_197(w_332_197, w_206_331, w_061_199);
  or2  I332_226(w_332_226, w_221_113, w_138_128);
  not1 I332_255(w_332_255, w_122_004);
  or2  I333_072(w_333_072, w_324_047, w_037_085);
  nand2 I333_074(w_333_074, w_165_004, w_004_346);
  not1 I333_091(w_333_091, w_219_011);
  or2  I333_179(w_333_179, w_043_143, w_318_342);
  nand2 I334_478(w_334_478, w_285_022, w_319_099);
  and2 I335_029(w_335_029, w_001_003, w_207_027);
  and2 I335_044(w_335_044, w_049_047, w_274_149);
  nand2 I335_066(w_335_066, w_049_329, w_272_020);
  and2 I335_091(w_335_091, w_149_003, w_162_010);
  not1 I335_121(w_335_121, w_263_026);
  or2  I335_209(w_335_209, w_150_082, w_142_131);
  or2  I336_060(w_336_060, w_230_053, w_155_102);
  not1 I336_091(w_336_091, w_130_087);
  not1 I336_289(w_336_289, w_146_245);
  not1 I336_307(w_336_307, w_034_076);
  not1 I337_030(w_337_030, w_092_156);
  not1 I337_118(w_337_118, w_273_143);
  and2 I337_195(w_337_195, w_036_016, w_159_073);
  not1 I337_215(w_337_215, w_210_032);
  or2  I338_026(w_338_026, w_189_029, w_095_051);
  or2  I338_063(w_338_063, w_084_055, w_087_188);
  or2  I338_069(w_338_069, w_284_265, w_061_032);
  and2 I338_278(w_338_278, w_241_021, w_255_057);
  not1 I338_330(w_338_330, w_308_024);
  and2 I338_356(w_338_358, w_333_074, w_338_357);
  nand2 I338_357(w_338_359, w_338_358, w_033_000);
  and2 I338_358(w_338_360, w_325_126, w_338_359);
  and2 I338_359(w_338_361, w_106_337, w_338_360);
  not1 I338_360(w_338_362, w_338_361);
  or2  I338_361(w_338_357, w_338_362, w_077_083);
  not1 I339_007(w_339_007, w_031_003);
  and2 I339_051(w_339_051, w_300_250, w_078_116);
  or2  I339_053(w_339_053, w_251_056, w_113_014);
  nand2 I339_177(w_339_177, w_309_065, w_135_027);
  nand2 I340_000(w_340_000, w_332_255, w_120_088);
  not1 I340_011(w_340_011, w_084_136);
  and2 I340_014(w_340_014, w_007_333, w_271_151);
  or2  I340_040(w_340_040, w_329_342, w_083_125);
  or2  I340_054(w_340_054, w_053_011, w_108_045);
  and2 I340_055(w_340_055, w_095_099, w_083_119);
  or2  I340_057(w_340_057, w_137_014, w_006_000);
  not1 I340_109(w_340_109, w_012_176);
  nand2 I341_000(w_341_000, w_250_044, w_166_021);
  or2  I342_008(w_342_008, w_242_346, w_253_140);
  nand2 I342_045(w_342_045, w_152_072, w_091_109);
  nand2 I342_047(w_342_047, w_323_046, w_340_055);
  and2 I342_126(w_342_126, w_081_025, w_077_162);
  and2 I342_127(w_342_127, w_304_065, w_000_439);
  nand2 I343_007(w_343_007, w_236_005, w_303_011);
  nand2 I343_037(w_343_037, w_219_300, w_208_126);
  nand2 I343_039(w_343_039, w_329_074, w_041_081);
  and2 I343_135(w_343_135, w_270_190, w_034_187);
  not1 I343_174(w_343_174, w_066_150);
  nand2 I343_228(w_343_228, w_228_066, w_041_164);
  and2 I343_266(w_343_266, w_131_127, w_336_091);
  and2 I344_173(w_344_173, w_231_066, w_031_067);
  not1 I344_199(w_344_199, w_167_302);
  not1 I344_457(w_344_457, w_137_045);
  and2 I345_011(w_345_011, w_271_338, w_248_133);
  not1 I345_135(w_345_135, w_139_187);
  nand2 I345_273(w_345_273, w_337_030, w_108_038);
  nand2 I345_274(w_345_274, w_312_123, w_130_068);
  not1 I346_050(w_346_050, w_131_081);
  nand2 I346_109(w_346_109, w_039_060, w_297_027);
  or2  I346_129(w_346_129, w_234_001, w_092_014);
  and2 I346_130(w_346_130, w_165_339, w_295_090);
  not1 I346_227(w_346_227, w_321_096);
  or2  I347_016(w_347_016, w_167_152, w_303_144);
  not1 I347_336(w_347_336, w_031_024);
  not1 I348_014(w_348_014, w_149_001);
  or2  I348_030(w_348_030, w_140_106, w_335_091);
  and2 I348_081(w_348_081, w_310_071, w_113_075);
  not1 I349_191(w_349_191, w_313_089);
  or2  I349_245(w_349_245, w_112_156, w_257_040);
  not1 I349_281(w_349_281, w_148_242);
  and2 I350_004(w_350_004, w_325_190, w_216_123);
  or2  I350_028(w_350_028, w_294_111, w_168_046);
  not1 I350_047(w_350_047, w_246_363);
  nand2 I350_238(w_350_238, w_177_212, w_016_380);
  nand2 I351_071(w_351_071, w_134_063, w_284_122);
  or2  I351_146(w_351_146, w_022_134, w_040_006);
  not1 I351_203(w_351_203, w_071_147);
  not1 I351_242(w_351_242, w_223_095);
  or2  I353_014(w_353_014, w_137_008, w_035_047);
  nand2 I353_076(w_353_076, w_204_066, w_305_057);
  nand2 I353_085(w_353_085, w_270_255, w_346_129);
  not1 I353_130(w_353_130, w_025_336);
  nand2 I354_003(w_354_003, w_166_181, w_061_160);
  not1 I354_039(w_354_039, w_107_047);
  and2 I354_041(w_354_041, w_313_074, w_267_389);
  and2 I354_079(w_354_079, w_307_123, w_319_064);
  and2 I355_015(w_355_015, w_170_038, w_345_274);
  not1 I355_017(w_355_017, w_038_049);
  and2 I355_028(w_355_028, w_220_054, w_127_172);
  nand2 I356_143(w_356_143, w_092_166, w_009_015);
  and2 I356_161(w_356_161, w_051_026, w_060_047);
  not1 I357_008(w_357_008, w_316_021);
  or2  I357_130(w_357_130, w_283_169, w_258_190);
  and2 I357_180(w_357_180, w_057_002, w_294_001);
  or2  I358_387(w_358_387, w_041_091, w_053_000);
  and2 I358_405(w_358_405, w_079_257, w_175_171);
  or2  I359_035(w_359_035, w_144_136, w_174_147);
  or2  I359_038(w_359_038, w_315_122, w_086_010);
  not1 I360_045(w_360_045, w_010_198);
  nand2 I360_064(w_360_064, w_323_057, w_229_092);
  or2  I360_083(w_360_083, w_152_032, w_062_002);
  not1 I360_088(w_360_088, w_116_100);
  nand2 I360_148(w_360_148, w_282_096, w_326_035);
  or2  I360_183(w_360_183, w_079_434, w_042_134);
  nand2 I361_066(w_361_066, w_120_021, w_287_308);
  or2  I361_099(w_361_099, w_254_101, w_359_038);
  and2 I362_046(w_362_046, w_283_026, w_320_219);
  or2  I362_069(w_362_069, w_066_169, w_010_283);
  not1 I363_010(w_363_010, w_008_081);
  nand2 I363_018(w_363_018, w_037_114, w_347_336);
  nand2 I363_068(w_363_068, w_155_101, w_038_030);
  and2 I363_072(w_363_072, w_013_195, w_171_276);
  not1 I363_094(w_363_094, w_065_121);
  or2  I363_100(w_363_100, w_036_034, w_179_138);
  and2 I364_037(w_364_037, w_210_176, w_121_001);
  not1 I364_083(w_364_083, w_239_236);
  nand2 I364_094(w_364_094, w_184_393, w_224_017);
  and2 I364_121(w_364_121, w_181_073, w_170_098);
  not1 I364_172(w_364_172, w_199_019);
  and2 I364_241(w_364_241, w_196_070, w_317_304);
  and2 I364_268(w_364_268, w_298_191, w_348_030);
  nand2 I365_028(w_365_028, w_044_018, w_192_221);
  not1 I365_042(w_365_042, w_210_226);
  not1 I365_077(w_365_077, w_070_055);
  and2 I365_141(w_365_141, w_013_208, w_088_435);
  or2  I366_026(w_366_026, w_215_234, w_044_158);
  or2  I366_124(w_366_124, w_121_070, w_043_129);
  nand2 I366_148(w_366_148, w_238_043, w_363_094);
  nand2 I366_183(w_366_183, w_129_000, w_059_346);
  and2 I366_193(w_366_193, w_191_075, w_260_074);
  not1 I366_206(w_366_206, w_008_195);
  and2 I367_049(w_367_049, w_297_016, w_059_191);
  or2  I367_165(w_367_165, w_042_016, w_096_154);
  or2  I367_393(w_367_393, w_250_029, w_035_035);
  or2  I368_097(w_368_097, w_165_111, w_354_041);
  or2  I368_099(w_368_099, w_097_097, w_212_052);
  nand2 I369_179(w_369_179, w_301_027, w_272_031);
  not1 I369_376(w_369_376, w_253_023);
  or2  I370_025(w_370_025, w_365_028, w_342_008);
  or2  I370_064(w_370_064, w_181_056, w_260_057);
  nand2 I370_123(w_370_123, w_302_029, w_085_027);
  and2 I370_137(w_370_137, w_199_018, w_193_039);
  or2  I371_122(w_371_122, w_014_043, w_093_034);
  not1 I371_325(w_371_325, w_136_002);
  and2 I372_024(w_372_024, w_172_018, w_290_019);
  and2 I372_062(w_372_062, w_264_085, w_127_404);
  or2  I372_070(w_372_070, w_024_105, w_161_207);
  and2 I372_146(w_372_148, w_372_147, w_315_242);
  or2  I372_147(w_372_149, w_372_148, w_205_047);
  and2 I372_148(w_372_150, w_372_149, w_316_057);
  nand2 I372_149(w_372_151, w_069_023, w_372_150);
  and2 I372_150(w_372_152, w_337_195, w_372_151);
  nand2 I372_151(w_372_153, w_372_152, w_309_115);
  nand2 I372_152(w_372_154, w_372_153, w_070_031);
  and2 I372_153(w_372_147, w_372_154, w_195_082);
  and2 I373_007(w_373_007, w_046_027, w_247_230);
  or2  I373_024(w_373_024, w_271_254, w_294_185);
  and2 I373_071(w_373_071, w_167_011, w_018_023);
  and2 I373_092(w_373_092, w_221_079, w_203_055);
  and2 I373_093(w_373_093, w_321_108, w_051_211);
  not1 I373_102(w_373_103, w_373_102);
  or2  I373_103(w_373_104, w_045_201, w_373_103);
  nand2 I373_104(w_373_105, w_373_104, w_103_012);
  or2  I373_105(w_373_106, w_127_033, w_373_105);
  nand2 I373_106(w_373_107, w_011_131, w_373_106);
  nand2 I373_107(w_373_102, w_373_107, w_188_109);
  or2  I374_002(w_374_002, w_139_030, w_178_121);
  and2 I374_034(w_374_034, w_323_033, w_339_051);
  not1 I374_035(w_374_035, w_056_071);
  and2 I374_110(w_374_110, w_263_053, w_267_222);
  and2 I375_169(w_375_169, w_018_162, w_176_396);
  nand2 I375_262(w_375_264, w_375_263, w_030_088);
  not1 I375_263(w_375_265, w_375_264);
  not1 I375_264(w_375_266, w_375_265);
  and2 I375_265(w_375_267, w_375_288, w_375_266);
  nand2 I375_266(w_375_268, w_182_024, w_375_267);
  or2  I375_267(w_375_269, w_375_268, w_316_044);
  nand2 I375_268(w_375_270, w_375_269, w_354_079);
  nand2 I375_269(w_375_271, w_375_270, w_370_064);
  not1 I375_270(w_375_272, w_375_271);
  not1 I375_271(w_375_263, w_375_272);
  or2  I375_272(w_375_277, w_139_188, w_375_276);
  not1 I375_273(w_375_278, w_375_277);
  and2 I375_274(w_375_279, w_224_053, w_375_278);
  not1 I375_275(w_375_280, w_375_279);
  and2 I375_276(w_375_281, w_028_188, w_375_280);
  and2 I375_277(w_375_282, w_003_061, w_375_281);
  or2  I375_278(w_375_283, w_375_282, w_313_119);
  nand2 I375_279(w_375_284, w_375_283, w_182_077);
  nand2 I375_280(w_375_285, w_374_035, w_375_284);
  or2  I375_281(w_375_286, w_009_033, w_375_285);
  not1 I375_282(w_375_276, w_375_267);
  and2 I375_283(w_375_288, w_073_117, w_375_286);
  or2  I376_092(w_376_092, w_012_365, w_142_078);
  or2  I376_151(w_376_151, w_268_018, w_340_054);
  and2 I377_008(w_377_008, w_163_000, w_272_003);
  not1 I377_053(w_377_053, w_150_156);
  nand2 I377_379(w_377_379, w_223_194, w_160_071);
  or2  I378_049(w_378_049, w_244_135, w_128_032);
  and2 I378_126(w_378_126, w_307_075, w_069_009);
  and2 I378_141(w_378_141, w_289_124, w_142_173);
  nand2 I378_179(w_378_179, w_007_164, w_219_246);
  nand2 I379_118(w_379_118, w_190_014, w_018_173);
  nand2 I380_152(w_380_152, w_120_004, w_224_012);
  nand2 I380_293(w_380_293, w_333_091, w_045_005);
  and2 I380_334(w_380_334, w_021_040, w_226_101);
  not1 I381_074(w_381_074, w_231_000);
  or2  I381_248(w_381_248, w_077_101, w_227_061);
  nand2 I381_443(w_381_443, w_214_029, w_220_358);
  or2  I382_002(w_382_002, w_221_046, w_373_093);
  nand2 I382_034(w_382_034, w_319_030, w_337_215);
  or2  I382_056(w_382_056, w_364_094, w_260_163);
  nand2 I383_159(w_383_159, w_279_071, w_089_031);
  and2 I384_042(w_384_042, w_111_020, w_111_024);
  or2  I384_057(w_384_057, w_240_206, w_231_041);
  and2 I384_072(w_384_072, w_161_153, w_093_365);
  and2 I385_013(w_385_013, w_061_337, w_300_121);
  and2 I385_014(w_385_014, w_059_440, w_196_211);
  nand2 I385_064(w_385_064, w_278_079, w_283_139);
  and2 I386_035(w_386_035, w_248_243, w_101_054);
  nand2 I386_178(w_386_178, w_280_063, w_280_008);
  and2 I386_290(w_386_290, w_171_227, w_360_045);
  and2 I387_024(w_387_024, w_287_423, w_179_084);
  nand2 I387_051(w_387_051, w_048_342, w_146_033);
  and2 I387_113(w_387_113, w_102_094, w_234_115);
  not1 I388_115(w_388_115, w_168_053);
  and2 I389_033(w_389_033, w_190_077, w_108_010);
  and2 I389_067(w_389_067, w_034_095, w_260_076);
  and2 I390_001(w_390_001, w_114_048, w_227_112);
  nand2 I390_052(w_390_052, w_059_341, w_377_379);
  and2 I392_137(w_392_137, w_160_075, w_342_126);
  or2  I392_288(w_392_288, w_221_099, w_335_066);
  nand2 I393_155(w_393_155, w_119_184, w_146_200);
  or2  I394_016(w_394_016, w_245_106, w_331_022);
  and2 I394_020(w_394_020, w_353_130, w_378_141);
  or2  I394_024(w_394_024, w_188_011, w_073_001);
  not1 I394_050(w_394_050, w_114_159);
  or2  I395_002(w_395_002, w_304_065, w_000_144);
  not1 I395_203(w_395_203, w_133_068);
  not1 I396_016(w_396_016, w_330_029);
  not1 I398_176(w_398_176, w_363_100);
  not1 I399_000(w_399_000, w_299_032);
  and2 I399_010(w_399_010, w_349_245, w_167_138);
  or2  I399_015(w_399_015, w_372_024, w_109_001);
  nand2 I399_028(w_399_028, w_334_478, w_168_054);
  nand2 I399_043(w_399_043, w_093_364, w_208_052);
  nand2 I399_049(w_399_049, w_357_130, w_072_014);
  nand2 I399_054(w_399_054, w_168_157, w_312_174);
  not1 I400_010(w_400_010, w_087_240);
  not1 I400_042(w_400_042, w_002_011);
  nand2 I400_047(w_400_047, w_006_000, w_093_004);
  and2 I400_075(w_400_075, w_263_040, w_372_062);
  and2 I400_084(w_400_084, w_065_032, w_252_092);
  not1 I400_091(w_400_091, w_370_025);
  and2 I401_091(w_401_091, w_384_072, w_208_037);
  or2  I401_410(w_401_410, w_363_072, w_213_177);
  not1 I402_009(w_402_009, w_251_113);
  not1 I402_035(w_402_035, w_157_242);
  nand2 I402_045(w_402_045, w_317_116, w_250_035);
  nand2 I403_036(w_403_036, w_028_130, w_172_041);
  and2 I404_279(w_404_279, w_014_008, w_366_183);
  not1 I404_377(w_404_377, w_009_129);
  not1 I405_041(w_405_041, w_266_314);
  and2 I405_167(w_405_167, w_093_346, w_307_002);
  or2  I405_178(w_405_178, w_164_020, w_171_268);
  or2  I407_015(w_407_015, w_312_171, w_176_380);
  nand2 I407_108(w_407_108, w_394_050, w_092_094);
  and2 I407_159(w_407_159, w_061_367, w_145_072);
  not1 I408_002(w_408_002, w_237_025);
  or2  I408_030(w_408_030, w_287_477, w_313_111);
  nand2 I408_171(w_408_171, w_257_168, w_226_310);
  not1 I408_216(w_408_216, w_002_011);
  nand2 I408_271(w_408_271, w_235_118, w_040_001);
  and2 I409_254(w_409_254, w_225_005, w_079_401);
  and2 I409_279(w_409_279, w_325_464, w_387_024);
  and2 I409_310(w_409_310, w_009_048, w_072_006);
  or2  I410_005(w_410_005, w_194_013, w_061_334);
  nand2 I410_075(w_410_075, w_105_057, w_252_279);
  not1 I411_149(w_411_149, w_343_007);
  nand2 I412_009(w_412_009, w_173_206, w_174_144);
  and2 I412_010(w_412_010, w_068_156, w_256_125);
  or2  I412_014(w_412_014, w_036_031, w_050_057);
  not1 I412_037(w_412_037, w_373_024);
  nand2 I413_022(w_413_022, w_018_158, w_274_192);
  or2  I413_029(w_413_029, w_307_062, w_024_194);
  not1 I413_052(w_413_052, w_263_194);
  or2  I413_064(w_413_064, w_158_001, w_294_037);
  or2  I414_028(w_414_028, w_180_133, w_086_084);
  or2  I415_029(w_415_029, w_215_228, w_219_290);
  and2 I415_041(w_415_041, w_060_064, w_328_215);
  and2 I415_054(w_415_054, w_314_142, w_259_102);
  not1 I416_296(w_416_296, w_254_037);
  or2  I416_319(w_416_319, w_343_039, w_349_281);
  and2 I416_450(w_416_450, w_272_029, w_039_151);
  not1 I417_006(w_417_006, w_289_089);
  and2 I417_038(w_417_038, w_178_104, w_211_075);
  nand2 I417_103(w_417_103, w_010_187, w_305_007);
  nand2 I417_133(w_417_133, w_381_248, w_147_066);
  or2  I418_069(w_418_069, w_079_219, w_343_037);
  not1 I418_107(w_418_107, w_400_047);
  not1 I418_144(w_418_144, w_333_179);
  and2 I419_064(w_419_064, w_283_224, w_240_041);
  or2  I420_044(w_420_044, w_215_102, w_139_043);
  or2  I420_081(w_420_081, w_272_010, w_131_169);
  nand2 I421_002(w_421_002, w_385_064, w_089_046);
  not1 I421_026(w_421_026, w_065_014);
  not1 I421_038(w_421_038, w_113_010);
  nand2 I421_047(w_421_047, w_321_056, w_308_027);
  not1 I421_048(w_421_048, w_415_054);
  or2  I421_063(w_421_063, w_091_152, w_202_032);
  nand2 I423_034(w_423_034, w_375_169, w_070_024);
  and2 I423_087(w_423_087, w_027_201, w_313_151);
  and2 I423_090(w_423_090, w_117_289, w_343_228);
  nand2 I423_096(w_423_096, w_293_134, w_033_028);
  or2  I424_100(w_424_100, w_360_064, w_138_223);
  and2 I425_154(w_425_154, w_188_105, w_033_051);
  nand2 I425_195(w_425_195, w_134_004, w_059_484);
  not1 I426_047(w_426_047, w_103_005);
  not1 I426_084(w_426_084, w_202_150);
  or2  I427_195(w_427_195, w_275_054, w_321_001);
  not1 I428_147(w_428_147, w_013_102);
  nand2 I428_176(w_428_176, w_004_054, w_173_062);
  not1 I428_202(w_428_202, w_289_118);
  nand2 I429_028(w_429_028, w_115_308, w_400_010);
  and2 I429_123(w_429_123, w_209_148, w_014_093);
  nand2 I429_342(w_429_342, w_402_009, w_029_012);
  or2  I430_100(w_430_100, w_183_036, w_034_031);
  or2  I430_237(w_430_237, w_092_171, w_208_022);
  nand2 I430_283(w_430_283, w_381_443, w_126_036);
  and2 I431_065(w_431_065, w_269_059, w_044_119);
  or2  I431_155(w_431_155, w_104_373, w_012_310);
  or2  I431_273(w_431_275, w_431_290, w_431_274);
  not1 I431_274(w_431_276, w_431_275);
  or2  I431_275(w_431_277, w_249_102, w_431_276);
  or2  I431_276(w_431_274, w_016_118, w_431_277);
  nand2 I431_277(w_431_282, w_246_078, w_431_281);
  not1 I431_278(w_431_283, w_431_282);
  and2 I431_279(w_431_284, w_431_283, w_172_094);
  and2 I431_280(w_431_285, w_431_284, w_393_155);
  and2 I431_281(w_431_286, w_431_285, w_115_185);
  or2  I431_282(w_431_287, w_013_160, w_431_286);
  not1 I431_283(w_431_288, w_431_287);
  not1 I431_284(w_431_281, w_431_275);
  and2 I431_285(w_431_290, w_079_235, w_431_288);
  not1 I432_071(w_432_071, w_104_374);
  not1 I432_131(w_432_131, w_360_148);
  nand2 I432_234(w_432_234, w_163_171, w_147_136);
  not1 I433_039(w_433_039, w_125_396);
  nand2 I433_297(w_433_297, w_242_105, w_065_210);
  or2  I434_098(w_434_098, w_257_048, w_203_235);
  or2  I434_174(w_434_174, w_316_014, w_096_283);
  nand2 I436_036(w_436_036, w_230_054, w_279_415);
  or2  I436_131(w_436_131, w_010_040, w_295_208);
  or2  I437_142(w_437_142, w_338_069, w_342_127);
  and2 I437_314(w_437_314, w_031_006, w_012_214);
  and2 I437_372(w_437_372, w_420_044, w_155_272);
  or2  I437_387(w_437_387, w_402_045, w_028_305);
  and2 I437_409(w_437_409, w_306_088, w_310_072);
  nand2 I438_037(w_438_037, w_270_111, w_364_121);
  not1 I439_040(w_439_040, w_409_279);
  or2  I439_186(w_439_186, w_330_154, w_373_092);
  nand2 I439_302(w_439_302, w_407_108, w_385_013);
  and2 I439_333(w_439_333, w_039_237, w_065_136);
  not1 I440_021(w_440_021, w_195_081);
  nand2 I440_090(w_440_090, w_259_131, w_322_030);
  and2 I441_005(w_441_005, w_060_226, w_111_001);
  or2  I441_048(w_441_048, w_367_393, w_338_278);
  and2 I441_160(w_441_160, w_363_010, w_382_056);
  nand2 I441_164(w_441_164, w_049_191, w_181_047);
  and2 I442_039(w_442_039, w_392_137, w_045_183);
  and2 I443_013(w_443_013, w_245_193, w_273_142);
  or2  I443_224(w_443_224, w_173_267, w_430_237);
  or2  I444_092(w_444_092, w_118_293, w_145_143);
  and2 I444_099(w_444_099, w_074_000, w_311_149);
  or2  I444_139(w_444_139, w_030_191, w_348_081);
  not1 I445_002(w_445_002, w_309_145);
  not1 I445_239(w_445_239, w_242_163);
  nand2 I445_354(w_445_354, w_282_037, w_256_072);
  nand2 I445_399(w_445_401, w_445_400, w_110_172);
  nand2 I445_400(w_445_402, w_445_401, w_445_416);
  or2  I445_401(w_445_403, w_292_099, w_445_402);
  and2 I445_402(w_445_404, w_298_112, w_445_403);
  nand2 I445_403(w_445_400, w_445_404, w_363_068);
  nand2 I445_404(w_445_409, w_178_104, w_445_408);
  or2  I445_405(w_445_410, w_445_409, w_185_122);
  not1 I445_406(w_445_411, w_445_410);
  nand2 I445_407(w_445_412, w_349_191, w_445_411);
  and2 I445_408(w_445_413, w_286_434, w_445_412);
  or2  I445_409(w_445_414, w_396_016, w_445_413);
  not1 I445_410(w_445_408, w_445_402);
  and2 I445_411(w_445_416, w_175_099, w_445_414);
  not1 I446_008(w_446_008, w_340_109);
  and2 I447_052(w_447_052, w_044_153, w_399_054);
  and2 I448_017(w_448_017, w_271_118, w_255_068);
  or2  I450_061(w_450_061, w_412_010, w_408_002);
  nand2 I450_294(w_450_294, w_032_045, w_256_134);
  not1 I452_024(w_452_024, w_178_049);
  and2 I452_134(w_452_134, w_428_176, w_329_287);
  not1 I453_014(w_453_014, w_012_014);
  or2  I453_051(w_453_051, w_260_063, w_147_019);
  not1 I453_349(w_453_349, w_272_009);
  and2 I454_080(w_454_080, w_383_159, w_338_026);
  not1 I454_088(w_454_088, w_008_061);
  nand2 I454_409(w_454_409, w_160_014, w_314_382);
  and2 I455_005(w_455_005, w_080_024, w_414_028);
  and2 I455_008(w_455_008, w_084_207, w_188_089);
  nand2 I455_023(w_455_023, w_298_031, w_163_147);
  nand2 I456_263(w_456_263, w_291_131, w_434_098);
  or2  I456_272(w_456_272, w_042_065, w_312_137);
  nand2 I456_397(w_456_397, w_076_009, w_182_026);
  and2 I458_002(w_458_002, w_395_002, w_202_411);
  nand2 I459_250(w_459_250, w_340_057, w_011_060);
  or2  I460_219(w_460_219, w_001_004, w_070_022);
  nand2 I461_097(w_461_097, w_140_005, w_029_028);
  nand2 I462_065(w_462_065, w_054_106, w_230_025);
  not1 I463_068(w_463_068, w_047_113);
  or2  I463_096(w_463_096, w_064_006, w_348_014);
  and2 I464_100(w_464_100, w_048_056, w_340_011);
  or2  I464_175(w_464_175, w_012_321, w_189_213);
  nand2 I465_019(w_465_019, w_207_204, w_082_032);
  or2  I467_079(w_467_079, w_115_095, w_351_242);
  not1 I467_208(w_467_208, w_122_021);
  and2 I467_415(w_467_415, w_194_058, w_156_168);
  nand2 I468_311(w_468_311, w_052_085, w_045_001);
  nand2 I468_341(w_468_341, w_314_369, w_344_457);
  not1 I468_377(w_468_377, w_188_048);
  and2 I469_026(w_469_026, w_128_058, w_249_033);
  or2  I469_317(w_469_317, w_304_188, w_354_039);
  not1 I469_331(w_469_331, w_107_041);
  not1 I471_034(w_471_034, w_380_152);
  nand2 I471_092(w_471_092, w_296_411, w_100_273);
  nand2 I472_120(w_472_120, w_326_040, w_275_088);
  not1 I473_338(w_473_338, w_442_039);
  not1 I474_062(w_474_062, w_249_031);
  nand2 I474_179(w_474_179, w_240_072, w_119_187);
  not1 I474_313(w_474_313, w_067_051);
  nand2 I475_091(w_475_091, w_341_000, w_322_007);
  and2 I475_104(w_475_104, w_051_045, w_411_149);
  nand2 I475_130(w_475_130, w_318_309, w_409_254);
  or2  I476_067(w_476_067, w_144_151, w_376_151);
  nand2 I476_251(w_476_253, w_476_252, w_222_218);
  not1 I476_252(w_476_254, w_476_253);
  nand2 I476_253(w_476_255, w_476_254, w_474_062);
  and2 I476_254(w_476_256, w_345_135, w_476_255);
  not1 I476_255(w_476_257, w_476_256);
  not1 I476_256(w_476_258, w_476_257);
  or2  I476_257(w_476_259, w_476_258, w_315_325);
  nand2 I476_258(w_476_260, w_016_225, w_476_259);
  and2 I476_259(w_476_252, w_206_030, w_476_260);
  not1 I477_036(w_477_036, w_025_194);
  or2  I477_047(w_477_047, w_075_081, w_033_001);
  and2 I478_218(w_478_218, w_030_049, w_013_073);
  or2  I478_276(w_478_276, w_208_076, w_248_029);
  nand2 I479_094(w_479_094, w_085_113, w_008_073);
  nand2 I480_000(w_480_000, w_026_206, w_286_002);
  or2  I480_002(w_480_002, w_458_002, w_430_100);
  nand2 I480_004(w_480_004, w_053_018, w_220_261);
  or2  I480_008(w_480_008, w_194_259, w_347_016);
  or2  I480_010(w_480_010, w_255_037, w_403_036);
  not1 I481_017(w_481_017, w_204_239);
  not1 I481_077(w_481_077, w_114_187);
  nand2 I482_000(w_482_000, w_332_197, w_312_222);
  not1 I482_001(w_482_001, w_027_138);
  and2 I482_008(w_482_008, w_381_074, w_218_163);
  and2 I483_015(w_483_015, w_327_163, w_434_174);
  not1 I483_041(w_483_041, w_247_254);
  not1 I484_029(w_484_029, w_225_167);
  and2 I484_091(w_484_093, w_484_092, w_012_081);
  nand2 I484_092(w_484_094, w_484_093, w_204_274);
  not1 I484_093(w_484_095, w_484_094);
  or2  I484_094(w_484_096, w_484_095, w_484_105);
  not1 I484_095(w_484_092, w_484_096);
  nand2 I484_096(w_484_101, w_484_100, w_417_133);
  not1 I484_097(w_484_102, w_484_101);
  not1 I484_098(w_484_103, w_484_102);
  not1 I484_099(w_484_100, w_484_096);
  and2 I484_100(w_484_105, w_421_002, w_484_103);
  nand2 I485_027(w_485_027, w_017_118, w_094_199);
  not1 I485_084(w_485_084, w_125_152);
  nand2 I486_007(w_486_007, w_309_073, w_462_065);
  and2 I487_030(w_487_030, w_146_064, w_080_011);
  or2  I487_053(w_487_053, w_190_066, w_119_040);
  and2 I487_054(w_487_054, w_298_024, w_052_023);
  and2 I487_064(w_487_064, w_338_330, w_387_113);
  not1 I487_076(w_487_078, w_487_077);
  nand2 I487_077(w_487_079, w_073_129, w_487_078);
  and2 I487_078(w_487_077, w_487_079, w_487_096);
  not1 I487_079(w_487_084, w_487_083);
  not1 I487_080(w_487_085, w_487_084);
  or2  I487_081(w_487_086, w_202_207, w_487_085);
  nand2 I487_082(w_487_087, w_003_054, w_487_086);
  not1 I487_083(w_487_088, w_487_087);
  nand2 I487_084(w_487_089, w_456_272, w_487_088);
  or2  I487_085(w_487_090, w_387_051, w_487_089);
  nand2 I487_086(w_487_091, w_358_405, w_487_090);
  nand2 I487_087(w_487_092, w_296_401, w_487_091);
  and2 I487_088(w_487_093, w_428_202, w_487_092);
  or2  I487_089(w_487_094, w_487_093, w_244_109);
  not1 I487_090(w_487_083, w_487_077);
  and2 I487_091(w_487_096, w_485_084, w_487_094);
  or2  I488_206(w_488_206, w_340_014, w_443_224);
  nand2 I489_322(w_489_324, w_489_323, w_346_109);
  or2  I489_323(w_489_325, w_489_344, w_489_324);
  nand2 I489_324(w_489_326, w_489_325, w_395_203);
  or2  I489_325(w_489_327, w_489_326, w_241_017);
  nand2 I489_326(w_489_328, w_426_047, w_489_327);
  not1 I489_327(w_489_329, w_489_328);
  or2  I489_328(w_489_330, w_489_329, w_201_196);
  and2 I489_329(w_489_331, w_489_330, w_183_077);
  nand2 I489_330(w_489_332, w_489_331, w_158_011);
  not1 I489_331(w_489_323, w_489_332);
  or2  I489_332(w_489_337, w_489_336, w_069_069);
  and2 I489_333(w_489_338, w_489_337, w_405_178);
  and2 I489_334(w_489_339, w_489_338, w_413_052);
  or2  I489_335(w_489_340, w_244_089, w_489_339);
  not1 I489_336(w_489_341, w_489_340);
  nand2 I489_337(w_489_342, w_489_341, w_423_096);
  not1 I489_338(w_489_336, w_489_325);
  and2 I489_339(w_489_344, w_187_131, w_489_342);
  nand2 I490_000(w_490_000, w_328_058, w_143_061);
  not1 I490_172(w_490_172, w_335_044);
  not1 I492_089(w_492_089, w_003_082);
  and2 I498_010(w_498_010, w_033_050, w_351_203);
  or2  I500_000(w_500_000, w_234_093, w_287_179);
  not1 I500_001(w_500_001, w_027_133);
  not1 I500_002(w_500_002, w_296_135);
  and2 I500_003(w_500_003, w_356_161, w_350_047);
  nand2 I500_004(w_500_004, w_265_003, w_240_180);
  and2 I500_005(w_500_005, w_071_036, w_054_038);
  nand2 I500_006(w_500_006, w_405_041, w_102_036);
  and2 I500_007(w_500_007, w_336_060, w_111_015);
  not1 I500_008(w_500_008, w_490_000);
  and2 I500_009(w_500_009, w_287_135, w_056_143);
  and2 I500_010(w_500_010, w_259_042, w_015_024);
  nand2 I500_011(w_500_011, w_108_024, w_400_084);
  or2  I500_012(w_500_012, w_306_287, w_020_024);
  not1 I500_013(w_500_013, w_123_067);
  nand2 I500_014(w_500_014, w_311_134, w_378_179);
  and2 I500_015(w_500_015, w_369_179, w_040_002);
  nand2 I500_016(w_500_016, w_096_151, w_167_037);
  or2  I500_017(w_500_017, w_035_038, w_413_064);
  and2 I500_018(w_500_018, w_165_174, w_029_223);
  or2  I500_019(w_500_019, w_402_035, w_404_377);
  or2  I500_020(w_500_020, w_319_081, w_231_049);
  nand2 I500_021(w_500_021, w_475_104, w_399_015);
  not1 I500_022(w_500_022, w_066_111);
  or2  I500_023(w_500_023, w_085_066, w_123_120);
  nand2 I500_024(w_500_024, w_388_115, w_487_053);
  or2  I500_025(w_500_025, w_369_376, w_103_005);
  nand2 I500_026(w_500_026, w_007_148, w_236_024);
  and2 I500_027(w_500_027, w_467_079, w_056_100);
  not1 I500_028(w_500_028, w_455_005);
  and2 I500_029(w_500_029, w_373_071, w_354_003);
  and2 I500_030(w_500_030, w_329_431, w_143_107);
  not1 I500_031(w_500_031, w_482_000);
  and2 I500_032(w_500_032, w_351_146, w_291_122);
  not1 I500_033(w_500_033, w_150_122);
  not1 I500_034(w_500_034, w_328_459);
  not1 I500_035(w_500_035, w_407_015);
  and2 I500_036(w_500_036, w_257_050, w_274_034);
  nand2 I500_037(w_500_037, w_399_000, w_153_001);
  or2  I500_038(w_500_038, w_436_036, w_286_039);
  and2 I500_039(w_500_039, w_408_171, w_172_168);
  not1 I500_040(w_500_040, w_146_168);
  and2 I500_041(w_500_041, w_269_043, w_292_087);
  or2  I500_042(w_500_042, w_051_095, w_301_161);
  or2  I500_043(w_500_043, w_075_047, w_464_100);
  nand2 I500_044(w_500_044, w_469_317, w_208_001);
  nand2 I500_045(w_500_045, w_346_130, w_124_106);
  and2 I500_046(w_500_046, w_148_012, w_374_002);
  or2  I500_047(w_500_047, w_338_063, w_200_130);
  nand2 I500_048(w_500_048, w_389_033, w_238_190);
  not1 I500_049(w_500_049, w_007_266);
  or2  I500_050(w_500_050, w_471_092, w_380_293);
  not1 I500_051(w_500_051, w_088_199);
  or2  I500_052(w_500_052, w_286_088, w_041_088);
  and2 I500_053(w_500_053, w_041_101, w_226_336);
  not1 I500_054(w_500_054, w_064_039);
  not1 I500_055(w_500_055, w_046_173);
  nand2 I500_056(w_500_056, w_079_133, w_069_108);
  or2  I500_057(w_500_057, w_187_053, w_316_046);
  and2 I500_058(w_500_058, w_109_000, w_188_047);
  nand2 I500_059(w_500_059, w_475_091, w_353_085);
  and2 I500_060(w_500_060, w_394_020, w_326_028);
  not1 I500_061(w_500_061, w_242_038);
  and2 I500_062(w_500_062, w_288_027, w_487_064);
  not1 I500_063(w_500_063, w_057_006);
  nand2 I500_064(w_500_064, w_096_017, w_024_228);
  or2  I500_065(w_500_065, w_485_027, w_150_146);
  not1 I500_066(w_500_066, w_125_246);
  nand2 I500_067(w_500_067, w_344_199, w_329_321);
  or2  I500_068(w_500_068, w_412_009, w_120_004);
  and2 I500_069(w_500_069, w_408_271, w_331_032);
  or2  I500_070(w_500_070, w_240_122, w_193_082);
  and2 I500_071(w_500_071, w_069_085, w_297_038);
  and2 I500_072(w_500_072, w_447_052, w_122_086);
  nand2 I500_073(w_500_073, w_057_060, w_350_238);
  not1 I500_074(w_500_074, w_227_150);
  or2  I500_075(w_500_075, w_199_006, w_373_007);
  nand2 I500_076(w_500_076, w_057_053, w_153_297);
  nand2 I500_077(w_500_077, w_346_227, w_047_267);
  and2 I500_078(w_500_078, w_344_173, w_296_144);
  not1 I500_079(w_500_079, w_418_144);
  or2  I500_080(w_500_080, w_327_041, w_431_065);
  nand2 I500_081(w_500_081, w_010_216, w_365_042);
  and2 I500_082(w_500_082, w_238_170, w_428_147);
  not1 I500_083(w_500_083, w_433_297);
  or2  I500_084(w_500_084, w_131_058, w_016_398);
  nand2 I500_085(w_500_085, w_213_071, w_335_209);
  or2  I500_086(w_500_086, w_105_129, w_230_017);
  nand2 I500_087(w_500_087, w_013_229, w_154_024);
  not1 I500_088(w_500_088, w_019_032);
  not1 I500_089(w_500_089, w_110_034);
  not1 I500_090(w_500_090, w_257_014);
  nand2 I500_091(w_500_091, w_054_048, w_170_190);
  and2 I500_092(w_500_092, w_420_081, w_417_038);
  or2  I500_093(w_500_093, w_126_009, w_374_110);
  and2 I500_094(w_500_094, w_307_129, w_089_305);
  or2  I500_095(w_500_095, w_465_019, w_453_051);
  or2  I500_096(w_500_096, w_415_029, w_452_024);
  not1 I500_097(w_500_097, w_343_135);
  not1 I500_098(w_500_098, w_366_193);
  not1 I500_099(w_500_099, w_286_054);
  and2 I500_100(w_500_100, w_130_146, w_258_046);
  not1 I500_101(w_500_101, w_366_124);
  or2  I500_102(w_500_102, w_293_011, w_162_007);
  nand2 I500_103(w_500_103, w_033_032, w_214_053);
  nand2 I500_104(w_500_104, w_374_034, w_323_000);
  not1 I500_105(w_500_105, w_106_262);
  and2 I500_106(w_500_106, w_079_328, w_382_034);
  and2 I500_107(w_500_107, w_365_141, w_071_193);
  nand2 I500_108(w_500_108, w_289_097, w_364_083);
  not1 I500_109(w_500_109, w_026_162);
  or2  I500_110(w_500_110, w_059_046, w_172_052);
  or2  I500_111(w_500_111, w_398_176, w_020_150);
  not1 I500_112(w_500_112, w_479_094);
  not1 I500_113(w_500_113, w_058_062);
  or2  I500_114(w_500_114, w_044_053, w_250_049);
  and2 I500_115(w_500_115, w_443_013, w_265_017);
  not1 I500_116(w_500_116, w_200_186);
  and2 I500_117(w_500_117, w_214_026, w_016_260);
  and2 I500_118(w_500_118, w_158_013, w_214_039);
  not1 I500_119(w_500_119, w_364_241);
  or2  I500_120(w_500_120, w_128_025, w_219_220);
  and2 I500_121(w_500_121, w_264_125, w_026_118);
  or2  I500_122(w_500_122, w_469_331, w_219_361);
  or2  I500_123(w_500_123, w_271_048, w_366_206);
  and2 I500_124(w_500_124, w_234_122, w_360_088);
  and2 I500_125(w_500_125, w_074_004, w_386_290);
  nand2 I500_126(w_500_126, w_195_080, w_211_135);
  not1 I500_127(w_500_127, w_487_030);
  and2 I500_128(w_500_128, w_366_148, w_421_063);
  and2 I500_129(w_500_129, w_140_049, w_093_264);
  or2  I500_130(w_500_130, w_459_250, w_141_193);
  and2 I500_131(w_500_131, w_353_014, w_404_279);
  and2 I500_132(w_500_132, w_290_069, w_483_015);
  nand2 I500_133(w_500_133, w_194_252, w_033_034);
  not1 I500_134(w_500_134, w_001_001);
  nand2 I500_135(w_500_135, w_423_087, w_467_415);
  and2 I500_136(w_500_136, w_060_179, w_437_372);
  or2  I500_137(w_500_137, w_078_081, w_130_106);
  nand2 I500_138(w_500_138, w_034_062, w_371_325);
  nand2 I500_139(w_500_139, w_206_162, w_174_253);
  not1 I500_140(w_500_140, w_208_004);
  or2  I500_141(w_500_141, w_061_039, w_036_204);
  not1 I500_142(w_500_142, w_355_028);
  nand2 I500_143(w_500_143, w_415_041, w_052_020);
  or2  I500_144(w_500_144, w_483_041, w_343_266);
  and2 I500_145(w_500_145, w_229_181, w_487_054);
  and2 I500_146(w_500_146, w_045_069, w_191_150);
  nand2 I500_147(w_500_147, w_399_049, w_440_021);
  and2 I500_148(w_500_148, w_328_297, w_307_183);
  or2  I500_149(w_500_149, w_274_017, w_184_178);
  not1 I500_150(w_500_150, w_249_052);
  nand2 I500_151(w_500_151, w_444_139, w_115_174);
  or2  I500_152(w_500_152, w_454_080, w_477_036);
  or2  I500_153(w_500_153, w_168_002, w_189_067);
  and2 I500_154(w_500_154, w_481_077, w_120_115);
  or2  I500_155(w_500_155, w_279_345, w_134_053);
  and2 I500_156(w_500_156, w_318_084, w_239_068);
  or2  I500_157(w_500_157, w_090_012, w_229_058);
  not1 I500_158(w_500_158, w_042_073);
  nand2 I500_159(w_500_159, w_372_070, w_268_040);
  nand2 I500_160(w_500_160, w_309_095, w_363_018);
  and2 I500_161(w_500_161, w_335_029, w_129_000);
  not1 I500_162(w_500_162, w_263_020);
  nand2 I500_163(w_500_163, w_081_001, w_390_001);
  not1 I500_164(w_500_164, w_480_002);
  nand2 I500_165(w_500_165, w_390_052, w_326_053);
  nand2 I500_166(w_500_166, w_198_323, w_440_090);
  not1 I500_167(w_500_167, w_101_254);
  or2  I500_168(w_500_168, w_096_150, w_445_002);
  nand2 I500_169(w_500_169, w_412_014, w_394_024);
  nand2 I500_170(w_500_170, w_328_241, w_093_329);
  nand2 I500_171(w_500_171, w_425_195, w_078_000);
  and2 I500_172(w_500_172, w_256_005, w_419_064);
  not1 I500_173(w_500_173, w_211_118);
  or2  I500_174(w_500_174, w_313_151, w_454_409);
  not1 I500_175(w_500_175, w_399_043);
  or2  I500_176(w_500_176, w_311_067, w_032_096);
  not1 I500_177(w_500_177, w_212_123);
  nand2 I500_178(w_500_178, w_041_132, w_492_089);
  not1 I500_179(w_500_179, w_012_337);
  nand2 I500_180(w_500_180, w_287_256, w_273_044);
  and2 I500_181(w_500_181, w_170_083, w_133_174);
  or2  I500_182(w_500_182, w_394_016, w_437_409);
  or2  I500_183(w_500_183, w_248_115, w_145_196);
  not1 I500_184(w_500_184, w_209_033);
  or2  I500_185(w_500_185, w_251_017, w_158_007);
  and2 I500_186(w_500_186, w_170_029, w_399_010);
  or2  I500_187(w_500_187, w_024_048, w_105_047);
  nand2 I500_188(w_500_188, w_090_221, w_168_151);
  or2  I500_189(w_500_189, w_105_246, w_014_206);
  nand2 I500_190(w_500_190, w_012_019, w_173_221);
  and2 I500_191(w_500_191, w_339_007, w_453_349);
  and2 I500_192(w_500_192, w_385_014, w_045_284);
  or2  I500_193(w_500_193, w_183_038, w_229_140);
  and2 I500_194(w_500_194, w_360_083, w_281_009);
  and2 I500_195(w_500_195, w_330_134, w_018_196);
  and2 I500_196(w_500_196, w_093_208, w_095_016);
  not1 I500_197(w_500_197, w_031_050);
  not1 I500_198(w_500_198, w_336_307);
  nand2 I500_199(w_500_199, w_222_030, w_020_171);
  and2 I500_200(w_500_200, w_055_019, w_441_048);
  nand2 I500_201(w_500_201, w_154_051, w_360_183);
  nand2 I500_202(w_500_202, w_042_169, w_125_239);
  not1 I500_203(w_500_203, w_071_299);
  or2  I500_204(w_500_204, w_190_081, w_340_000);
  and2 I500_205(w_500_205, w_028_159, w_163_250);
  or2  I500_206(w_500_206, w_035_005, w_401_091);
  and2 I500_207(w_500_207, w_195_016, w_412_037);
  not1 I500_208(w_500_208, w_272_024);
  or2  I500_209(w_500_209, w_167_053, w_206_063);
  nand2 I500_210(w_500_210, w_277_005, w_076_077);
  nand2 I500_211(w_500_211, w_416_319, w_327_176);
  not1 I500_212(w_500_212, w_342_047);
  and2 I500_213(w_500_213, w_377_008, w_421_048);
  or2  I500_214(w_500_214, w_468_311, w_105_317);
  or2  I500_215(w_500_215, w_377_053, w_218_396);
  nand2 I500_216(w_500_216, w_425_154, w_226_202);
  and2 I500_217(w_500_217, w_303_178, w_351_071);
  or2  I500_218(w_500_218, w_030_016, w_024_071);
  and2 I500_219(w_500_219, w_044_101, w_276_117);
  not1 I500_220(w_500_220, w_117_434);
  or2  I500_221(w_500_221, w_074_001, w_223_099);
  or2  I500_222(w_500_222, w_441_005, w_116_218);
  nand2 I500_223(w_500_223, w_194_273, w_067_035);
  nand2 I500_224(w_500_224, w_418_069, w_340_040);
  or2  I500_225(w_500_225, w_364_172, w_205_023);
  or2  I500_226(w_500_226, w_482_001, w_047_015);
  and2 I500_227(w_500_227, w_133_026, w_467_208);
  not1 I500_228(w_500_228, w_124_001);
  not1 I500_229(w_500_229, w_092_033);
  or2  I500_230(w_500_230, w_287_000, w_304_136);
  and2 I500_231(w_500_231, w_074_003, w_332_226);
  nand2 I500_232(w_500_232, w_049_250, w_052_071);
  and2 I500_233(w_500_233, w_386_035, w_423_090);
  nand2 I500_234(w_500_234, w_408_216, w_367_049);
  not1 I500_235(w_500_235, w_343_174);
  and2 I500_236(w_500_236, w_288_190, w_370_137);
  nand2 I500_237(w_500_237, w_174_063, w_027_101);
  or2  I500_238(w_500_238, w_359_035, w_320_260);
  not1 I500_239(w_500_239, w_224_000);
  not1 I500_240(w_500_240, w_463_068);
  or2  I500_241(w_500_241, w_153_209, w_342_045);
  and2 I500_242(w_500_242, w_310_226, w_271_280);
  nand2 I500_243(w_500_243, w_059_322, w_473_338);
  or2  I500_244(w_500_244, w_000_402, w_236_068);
  nand2 I500_245(w_500_245, w_448_017, w_399_028);
  not1 I500_246(w_500_246, w_475_130);
  and2 I500_247(w_500_247, w_438_037, w_450_061);
  or2  I500_248(w_500_248, w_144_016, w_077_201);
  nand2 I500_249(w_500_249, w_200_235, w_091_260);
  or2  I500_250(w_500_250, w_416_450, w_119_122);
  and2 I500_251(w_500_251, w_355_017, w_431_155);
  not1 I500_252(w_500_252, w_330_364);
  and2 I500_253(w_500_253, w_306_004, w_137_035);
  not1 I500_254(w_500_254, w_439_040);
  nand2 I500_255(w_500_255, w_083_188, w_364_037);
  and2 I500_256(w_500_256, w_065_124, w_339_177);
  not1 I500_257(w_500_257, w_107_057);
  or2  I500_258(w_500_258, w_024_031, w_212_031);
  nand2 I500_259(w_500_259, w_368_099, w_446_008);
  and2 I500_260(w_500_260, w_104_430, w_005_200);
  or2  I500_261(w_500_261, w_444_092, w_004_027);
  or2  I500_262(w_500_262, w_221_064, w_249_029);
  or2  I500_263(w_500_263, w_088_315, w_427_195);
  not1 I500_264(w_500_264, w_432_071);
  not1 I500_265(w_500_265, w_144_124);
  not1 I500_266(w_500_266, w_364_268);
  and2 I500_267(w_500_267, w_096_136, w_144_186);
  or2  I500_268(w_500_268, w_196_096, w_085_036);
  and2 I500_269(w_500_269, w_112_142, w_025_029);
  nand2 I500_270(w_500_270, w_163_070, w_331_042);
  or2  I500_271(w_500_271, w_026_125, w_281_010);
  nand2 I500_272(w_500_272, w_277_015, w_197_142);
  nand2 I500_273(w_500_273, w_089_090, w_024_085);
  or2  I500_274(w_500_274, w_165_282, w_417_103);
  nand2 I500_275(w_500_275, w_222_067, w_065_021);
  and2 I500_276(w_500_276, w_456_263, w_018_287);
  or2  I500_277(w_500_277, w_367_165, w_070_000);
  nand2 I500_278(w_500_278, w_174_278, w_234_099);
  and2 I500_279(w_500_279, w_474_313, w_362_046);
  not1 I500_280(w_500_280, w_184_015);
  and2 I500_281(w_500_281, w_453_014, w_455_023);
  not1 I500_282(w_500_282, w_020_088);
  not1 I500_283(w_500_283, w_328_038);
  or2  I500_284(w_500_284, w_115_131, w_224_001);
  not1 I500_285(w_500_285, w_225_248);
  and2 I500_286(w_500_286, w_355_015, w_303_127);
  or2  I500_287(w_500_287, w_468_341, w_159_072);
  or2  I500_288(w_500_288, w_026_251, w_331_017);
  nand2 I500_289(w_500_289, w_358_387, w_079_133);
  or2  I500_290(w_500_290, w_408_171, w_378_126);
  nand2 I500_291(w_500_291, w_455_008, w_357_180);
  or2  I500_292(w_500_292, w_437_387, w_444_099);
  not1 I500_293(w_500_293, w_253_048);
  nand2 I500_294(w_500_294, w_264_064, w_437_142);
  nand2 I500_295(w_500_295, w_268_139, w_238_126);
  not1 I500_296(w_500_296, w_170_112);
  and2 I500_297(w_500_297, w_430_283, w_482_008);
  not1 I500_298(w_500_298, w_437_314);
  nand2 I500_299(w_500_299, w_469_026, w_436_131);
  nand2 I500_300(w_500_300, w_177_222, w_120_043);
  not1 I500_301(w_500_301, w_236_018);
  nand2 I500_302(w_500_302, w_378_049, w_339_053);
  and2 I500_303(w_500_303, w_317_248, w_310_184);
  and2 I500_304(w_500_304, w_240_213, w_335_121);
  nand2 I500_305(w_500_305, w_124_211, w_003_094);
  not1 I500_306(w_500_306, w_439_302);
  or2  I500_307(w_500_307, w_468_377, w_325_206);
  nand2 I500_308(w_500_308, w_061_224, w_230_043);
  not1 I500_309(w_500_309, w_421_026);
  not1 I500_310(w_500_310, w_238_262);
  and2 I500_311(w_500_311, w_168_115, w_168_047);
  not1 I500_312(w_500_312, w_065_010);
  not1 I500_313(w_500_313, w_129_000);
  and2 I500_314(w_500_314, w_115_031, w_027_321);
  nand2 I500_315(w_500_315, w_256_011, w_058_000);
  and2 I500_316(w_500_316, w_134_022, w_204_260);
  not1 I500_317(w_500_317, w_366_026);
  and2 I500_318(w_500_318, w_480_010, w_028_049);
  not1 I500_319(w_500_319, w_261_115);
  and2 I500_320(w_500_320, w_350_028, w_021_105);
  and2 I500_321(w_500_321, w_488_206, w_279_309);
  and2 I500_322(w_500_322, w_035_080, w_382_002);
  and2 I500_323(w_500_323, w_016_151, w_424_100);
  or2  I500_324(w_500_324, w_142_303, w_282_122);
  not1 I500_325(w_500_325, w_310_070);
  and2 I500_326(w_500_326, w_072_064, w_272_022);
  nand2 I500_327(w_500_327, w_145_215, w_452_134);
  and2 I500_328(w_500_328, w_083_003, w_012_119);
  nand2 I500_329(w_500_329, w_246_273, w_175_262);
  or2  I500_330(w_500_330, w_099_088, w_198_093);
  nand2 I500_331(w_500_331, w_480_008, w_305_054);
  not1 I500_332(w_500_332, w_389_067);
  or2  I500_333(w_500_333, w_162_001, w_361_099);
  and2 I500_334(w_500_334, w_165_293, w_096_248);
  or2  I500_335(w_500_335, w_460_219, w_192_206);
  or2  I500_336(w_500_336, w_368_097, w_270_054);
  and2 I500_337(w_500_337, w_320_108, w_259_153);
  or2  I500_338(w_500_338, w_416_296, w_471_034);
  nand2 I500_339(w_500_339, w_132_054, w_056_151);
  nand2 I500_340(w_500_340, w_464_175, w_273_071);
  nand2 I500_341(w_500_341, w_362_069, w_182_100);
  and2 I500_342(w_500_342, w_175_274, w_105_297);
  not1 I500_343(w_500_343, w_169_217);
  nand2 I500_344(w_500_344, w_429_123, w_192_086);
  nand2 I500_345(w_500_345, w_163_003, w_486_007);
  nand2 I500_346(w_500_346, w_042_054, w_303_162);
  nand2 I500_347(w_500_347, w_076_029, w_318_290);
  or2  I500_348(w_500_348, w_001_000, w_429_028);
  nand2 I500_349(w_500_349, w_386_178, w_269_055);
  and2 I500_350(w_500_350, w_480_004, w_271_172);
  not1 I500_351(w_500_351, w_042_187);
  or2  I500_352(w_500_352, w_380_334, w_361_066);
  nand2 I500_353(w_500_353, w_164_132, w_239_092);
  and2 I500_354(w_500_354, w_057_016, w_401_410);
  not1 I500_355(w_500_355, w_182_087);
  or2  I500_356(w_500_356, w_068_155, w_022_149);
  or2  I500_357(w_500_357, w_002_004, w_240_026);
  not1 I500_358(w_500_358, w_282_065);
  nand2 I500_359(w_500_359, w_014_252, w_392_288);
  nand2 I500_360(w_500_360, w_408_030, w_022_000);
  and2 I500_361(w_500_361, w_432_234, w_429_342);
  or2  I500_362(w_500_362, w_463_096, w_418_107);
  not1 I500_363(w_500_363, w_441_164);
  nand2 I500_364(w_500_364, w_295_171, w_311_174);
  or2  I500_365(w_500_365, w_445_239, w_048_071);
  nand2 I500_366(w_500_366, w_293_099, w_275_053);
  and2 I500_367(w_500_367, w_149_000, w_048_081);
  and2 I500_368(w_500_368, w_478_276, w_305_085);
  or2  I500_369(w_500_369, w_224_045, w_216_017);
  and2 I500_370(w_500_370, w_139_164, w_207_303);
  not1 I500_371(w_500_371, w_224_038);
  not1 I500_372(w_500_372, w_272_024);
  or2  I500_373(w_500_373, w_417_006, w_400_091);
  nand2 I500_374(w_500_374, w_050_172, w_432_131);
  or2  I500_375(w_500_375, w_410_075, w_175_203);
  or2  I500_376(w_500_376, w_251_124, w_089_120);
  and2 I500_377(w_500_377, w_228_284, w_123_012);
  nand2 I500_378(w_500_378, w_199_018, w_257_052);
  and2 I500_379(w_500_379, w_030_041, w_055_083);
  and2 I500_380(w_500_380, w_439_333, w_293_037);
  and2 I500_381(w_500_381, w_163_133, w_076_069);
  and2 I500_382(w_500_382, w_097_193, w_421_038);
  or2  I500_383(w_500_383, w_337_118, w_197_083);
  not1 I500_384(w_500_384, w_172_012);
  not1 I500_385(w_500_385, w_281_016);
  not1 I500_386(w_500_386, w_312_199);
  or2  I500_387(w_500_387, w_095_037, w_376_092);
  and2 I500_388(w_500_388, w_099_244, w_303_084);
  and2 I500_389(w_500_389, w_345_273, w_269_038);
  not1 I500_390(w_500_390, w_159_199);
  nand2 I500_391(w_500_391, w_278_118, w_048_280);
  or2  I500_392(w_500_392, w_413_029, w_054_101);
  and2 I500_393(w_500_393, w_218_031, w_085_060);
  not1 I500_394(w_500_394, w_314_093);
  not1 I500_395(w_500_395, w_413_022);
  or2  I500_396(w_500_396, w_498_010, w_370_123);
  and2 I500_397(w_500_397, w_008_169, w_291_015);
  and2 I500_398(w_500_398, w_421_047, w_101_201);
  and2 I500_399(w_500_399, w_014_053, w_135_115);
  nand2 I500_400(w_500_400, w_353_076, w_405_167);
  or2  I500_401(w_500_401, w_219_260, w_099_181);
  not1 I500_402(w_500_402, w_124_088);
  or2  I500_403(w_500_403, w_346_050, w_445_354);
  not1 I500_404(w_500_404, w_088_061);
  nand2 I500_405(w_500_405, w_010_368, w_484_029);
  or2  I500_406(w_500_406, w_350_004, w_084_114);
  not1 I500_407(w_500_407, w_289_120);
  nand2 I500_408(w_500_408, w_456_397, w_326_069);
  and2 I500_409(w_500_409, w_163_371, w_472_120);
  and2 I500_410(w_500_410, w_318_159, w_481_017);
  or2  I500_411(w_500_411, w_070_085, w_020_080);
  not1 I500_412(w_500_412, w_356_143);
  nand2 I500_413(w_500_413, w_206_035, w_191_024);
  or2  I500_414(w_500_414, w_332_014, w_336_289);
  not1 I500_415(w_500_415, w_015_074);
  not1 I500_416(w_500_416, w_030_081);
  nand2 I500_417(w_500_417, w_379_118, w_081_026);
  nand2 I500_418(w_500_418, w_106_232, w_021_079);
  and2 I500_419(w_500_419, w_101_002, w_461_097);
  and2 I500_420(w_500_420, w_167_157, w_147_191);
  and2 I500_421(w_500_421, w_480_000, w_245_121);
  not1 I500_422(w_500_422, w_260_000);
  and2 I500_423(w_500_423, w_142_116, w_175_373);
  not1 I500_424(w_500_424, w_109_000);
  not1 I500_425(w_500_425, w_215_054);
  nand2 I500_426(w_500_426, w_258_022, w_161_171);
  or2  I500_427(w_500_427, w_110_194, w_081_073);
  and2 I500_428(w_500_428, w_124_002, w_248_360);
  nand2 I500_429(w_500_429, w_221_050, w_203_038);
  nand2 I500_430(w_500_430, w_345_011, w_478_218);
  nand2 I500_431(w_500_431, w_439_186, w_145_006);
  not1 I500_432(w_500_432, w_204_117);
  nand2 I500_433(w_500_433, w_365_077, w_400_042);
  or2  I500_434(w_500_434, w_333_072, w_409_310);
  nand2 I500_435(w_500_435, w_009_170, w_202_230);
  or2  I500_436(w_500_436, w_257_214, w_160_102);
  nand2 I500_437(w_500_437, w_490_172, w_318_049);
  nand2 I500_438(w_500_438, w_315_288, w_245_019);
  or2  I500_439(w_500_439, w_232_075, w_482_008);
  and2 I500_440(w_500_440, w_476_067, w_329_237);
  and2 I500_441(w_500_441, w_292_106, w_151_034);
  or2  I500_442(w_500_442, w_212_037, w_316_224);
  or2  I500_443(w_500_443, w_175_214, w_230_013);
  and2 I500_444(w_500_444, w_441_160, w_285_018);
  nand2 I500_445(w_500_445, w_190_025, w_268_025);
  and2 I500_446(w_500_446, w_185_031, w_426_084);
  not1 I500_447(w_500_447, w_407_159);
  or2  I500_448(w_500_448, w_410_005, w_371_122);
  or2  I500_449(w_500_449, w_187_032, w_314_214);
  and2 I500_450(w_500_450, w_044_059, w_261_083);
  nand2 I500_451(w_500_451, w_046_024, w_454_088);
  nand2 I500_452(w_500_452, w_075_113, w_051_260);
  not1 I500_453(w_500_453, w_477_047);
  or2  I500_454(w_500_454, w_384_042, w_450_294);
  nand2 I500_455(w_500_455, w_173_134, w_400_075);
  not1 I500_456(w_500_456, w_066_074);
  nand2 I500_457(w_500_457, w_463_096, w_140_300);
  and2 I500_458(w_500_458, w_186_024, w_011_126);
  nand2 I500_459(w_500_459, w_086_092, w_170_198);
  not1 I500_460(w_500_460, w_148_324);
  nand2 I500_461(w_500_461, w_384_057, w_474_179);
  or2  I500_462(w_500_462, w_147_063, w_357_008);
  not1 I500_463(w_500_463, w_423_034);
  or2  I500_464(w_500_464, w_238_272, w_433_039);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_300, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_328, w_000_330, w_000_331, w_000_332, w_000_335, w_000_336, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_356, w_000_358, w_000_359, w_000_360, w_000_363, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_420, w_000_422, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_431, w_000_433, w_000_434, w_000_437, w_000_439, w_000_440, w_000_444, w_000_445, w_000_447, w_000_448, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_457, w_000_458, w_000_462, w_000_463, w_000_468, w_000_474, w_000_490, w_500_000, w_500_001, w_500_002, w_500_003, w_500_004, w_500_005, w_500_006, w_500_007, w_500_008, w_500_009, w_500_010, w_500_011, w_500_012, w_500_013, w_500_014, w_500_015, w_500_016, w_500_017, w_500_018, w_500_019, w_500_020, w_500_021, w_500_022, w_500_023, w_500_024, w_500_025, w_500_026, w_500_027, w_500_028, w_500_029, w_500_030, w_500_031, w_500_032, w_500_033, w_500_034, w_500_035, w_500_036, w_500_037, w_500_038, w_500_039, w_500_040, w_500_041, w_500_042, w_500_043, w_500_044, w_500_045, w_500_046, w_500_047, w_500_048, w_500_049, w_500_050, w_500_051, w_500_052, w_500_053, w_500_054, w_500_055, w_500_056, w_500_057, w_500_058, w_500_059, w_500_060, w_500_061, w_500_062, w_500_063, w_500_064, w_500_065, w_500_066, w_500_067, w_500_068, w_500_069, w_500_070, w_500_071, w_500_072, w_500_073, w_500_074, w_500_075, w_500_076, w_500_077, w_500_078, w_500_079, w_500_080, w_500_081, w_500_082, w_500_083, w_500_084, w_500_085, w_500_086, w_500_087, w_500_088, w_500_089, w_500_090, w_500_091, w_500_092, w_500_093, w_500_094, w_500_095, w_500_096, w_500_097, w_500_098, w_500_099, w_500_100, w_500_101, w_500_102, w_500_103, w_500_104, w_500_105, w_500_106, w_500_107, w_500_108, w_500_109, w_500_110, w_500_111, w_500_112, w_500_113, w_500_114, w_500_115, w_500_116, w_500_117, w_500_118, w_500_119, w_500_120, w_500_121, w_500_122, w_500_123, w_500_124, w_500_125, w_500_126, w_500_127, w_500_128, w_500_129, w_500_130, w_500_131, w_500_132, w_500_133, w_500_134, w_500_135, w_500_136, w_500_137, w_500_138, w_500_139, w_500_140, w_500_141, w_500_142, w_500_143, w_500_144, w_500_145, w_500_146, w_500_147, w_500_148, w_500_149, w_500_150, w_500_151, w_500_152, w_500_153, w_500_154, w_500_155, w_500_156, w_500_157, w_500_158, w_500_159, w_500_160, w_500_161, w_500_162, w_500_163, w_500_164, w_500_165, w_500_166, w_500_167, w_500_168, w_500_169, w_500_170, w_500_171, w_500_172, w_500_173, w_500_174, w_500_175, w_500_176, w_500_177, w_500_178, w_500_179, w_500_180, w_500_181, w_500_182, w_500_183, w_500_184, w_500_185, w_500_186, w_500_187, w_500_188, w_500_189, w_500_190, w_500_191, w_500_192, w_500_193, w_500_194, w_500_195, w_500_196, w_500_197, w_500_198, w_500_199, w_500_200, w_500_201, w_500_202, w_500_203, w_500_204, w_500_205, w_500_206, w_500_207, w_500_208, w_500_209, w_500_210, w_500_211, w_500_212, w_500_213, w_500_214, w_500_215, w_500_216, w_500_217, w_500_218, w_500_219, w_500_220, w_500_221, w_500_222, w_500_223, w_500_224, w_500_225, w_500_226, w_500_227, w_500_228, w_500_229, w_500_230, w_500_231, w_500_232, w_500_233, w_500_234, w_500_235, w_500_236, w_500_237, w_500_238, w_500_239, w_500_240, w_500_241, w_500_242, w_500_243, w_500_244, w_500_245, w_500_246, w_500_247, w_500_248, w_500_249, w_500_250, w_500_251, w_500_252, w_500_253, w_500_254, w_500_255, w_500_256, w_500_257, w_500_258, w_500_259, w_500_260, w_500_261, w_500_262, w_500_263, w_500_264, w_500_265, w_500_266, w_500_267, w_500_268, w_500_269, w_500_270, w_500_271, w_500_272, w_500_273, w_500_274, w_500_275, w_500_276, w_500_277, w_500_278, w_500_279, w_500_280, w_500_281, w_500_282, w_500_283, w_500_284, w_500_285, w_500_286, w_500_287, w_500_288, w_500_289, w_500_290, w_500_291, w_500_292, w_500_293, w_500_294, w_500_295, w_500_296, w_500_297, w_500_298, w_500_299, w_500_300, w_500_301, w_500_302, w_500_303, w_500_304, w_500_305, w_500_306, w_500_307, w_500_308, w_500_309, w_500_310, w_500_311, w_500_312, w_500_313, w_500_314, w_500_315, w_500_316, w_500_317, w_500_318, w_500_319, w_500_320, w_500_321, w_500_322, w_500_323, w_500_324, w_500_325, w_500_326, w_500_327, w_500_328, w_500_329, w_500_330, w_500_331, w_500_332, w_500_333, w_500_334, w_500_335, w_500_336, w_500_337, w_500_338, w_500_339, w_500_340, w_500_341, w_500_342, w_500_343, w_500_344, w_500_345, w_500_346, w_500_347, w_500_348, w_500_349, w_500_350, w_500_351, w_500_352, w_500_353, w_500_354, w_500_355, w_500_356, w_500_357, w_500_358, w_500_359, w_500_360, w_500_361, w_500_362, w_500_363, w_500_364, w_500_365, w_500_366, w_500_367, w_500_368, w_500_369, w_500_370, w_500_371, w_500_372, w_500_373, w_500_374, w_500_375, w_500_376, w_500_377, w_500_378, w_500_379, w_500_380, w_500_381, w_500_382, w_500_383, w_500_384, w_500_385, w_500_386, w_500_387, w_500_388, w_500_389, w_500_390, w_500_391, w_500_392, w_500_393, w_500_394, w_500_395, w_500_396, w_500_397, w_500_398, w_500_399, w_500_400, w_500_401, w_500_402, w_500_403, w_500_404, w_500_405, w_500_406, w_500_407, w_500_408, w_500_409, w_500_410, w_500_411, w_500_412, w_500_413, w_500_414, w_500_415, w_500_416, w_500_417, w_500_418, w_500_419, w_500_420, w_500_421, w_500_422, w_500_423, w_500_424, w_500_425, w_500_426, w_500_427, w_500_428, w_500_429, w_500_430, w_500_431, w_500_432, w_500_433, w_500_434, w_500_435, w_500_436, w_500_437, w_500_438, w_500_439, w_500_440, w_500_441, w_500_442, w_500_443, w_500_444, w_500_445, w_500_446, w_500_447, w_500_448, w_500_449, w_500_450, w_500_451, w_500_452, w_500_453, w_500_454, w_500_455, w_500_456, w_500_457, w_500_458, w_500_459, w_500_460, w_500_461, w_500_462, w_500_463, w_500_464 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_300, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_328, w_000_330, w_000_331, w_000_332, w_000_335, w_000_336, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_356, w_000_358, w_000_359, w_000_360, w_000_363, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_420, w_000_422, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_431, w_000_433, w_000_434, w_000_437, w_000_439, w_000_440, w_000_444, w_000_445, w_000_447, w_000_448, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_457, w_000_458, w_000_462, w_000_463, w_000_468, w_000_474, w_000_490, w_500_000, w_500_001, w_500_002, w_500_003, w_500_004, w_500_005, w_500_006, w_500_007, w_500_008, w_500_009, w_500_010, w_500_011, w_500_012, w_500_013, w_500_014, w_500_015, w_500_016, w_500_017, w_500_018, w_500_019, w_500_020, w_500_021, w_500_022, w_500_023, w_500_024, w_500_025, w_500_026, w_500_027, w_500_028, w_500_029, w_500_030, w_500_031, w_500_032, w_500_033, w_500_034, w_500_035, w_500_036, w_500_037, w_500_038, w_500_039, w_500_040, w_500_041, w_500_042, w_500_043, w_500_044, w_500_045, w_500_046, w_500_047, w_500_048, w_500_049, w_500_050, w_500_051, w_500_052, w_500_053, w_500_054, w_500_055, w_500_056, w_500_057, w_500_058, w_500_059, w_500_060, w_500_061, w_500_062, w_500_063, w_500_064, w_500_065, w_500_066, w_500_067, w_500_068, w_500_069, w_500_070, w_500_071, w_500_072, w_500_073, w_500_074, w_500_075, w_500_076, w_500_077, w_500_078, w_500_079, w_500_080, w_500_081, w_500_082, w_500_083, w_500_084, w_500_085, w_500_086, w_500_087, w_500_088, w_500_089, w_500_090, w_500_091, w_500_092, w_500_093, w_500_094, w_500_095, w_500_096, w_500_097, w_500_098, w_500_099, w_500_100, w_500_101, w_500_102, w_500_103, w_500_104, w_500_105, w_500_106, w_500_107, w_500_108, w_500_109, w_500_110, w_500_111, w_500_112, w_500_113, w_500_114, w_500_115, w_500_116, w_500_117, w_500_118, w_500_119, w_500_120, w_500_121, w_500_122, w_500_123, w_500_124, w_500_125, w_500_126, w_500_127, w_500_128, w_500_129, w_500_130, w_500_131, w_500_132, w_500_133, w_500_134, w_500_135, w_500_136, w_500_137, w_500_138, w_500_139, w_500_140, w_500_141, w_500_142, w_500_143, w_500_144, w_500_145, w_500_146, w_500_147, w_500_148, w_500_149, w_500_150, w_500_151, w_500_152, w_500_153, w_500_154, w_500_155, w_500_156, w_500_157, w_500_158, w_500_159, w_500_160, w_500_161, w_500_162, w_500_163, w_500_164, w_500_165, w_500_166, w_500_167, w_500_168, w_500_169, w_500_170, w_500_171, w_500_172, w_500_173, w_500_174, w_500_175, w_500_176, w_500_177, w_500_178, w_500_179, w_500_180, w_500_181, w_500_182, w_500_183, w_500_184, w_500_185, w_500_186, w_500_187, w_500_188, w_500_189, w_500_190, w_500_191, w_500_192, w_500_193, w_500_194, w_500_195, w_500_196, w_500_197, w_500_198, w_500_199, w_500_200, w_500_201, w_500_202, w_500_203, w_500_204, w_500_205, w_500_206, w_500_207, w_500_208, w_500_209, w_500_210, w_500_211, w_500_212, w_500_213, w_500_214, w_500_215, w_500_216, w_500_217, w_500_218, w_500_219, w_500_220, w_500_221, w_500_222, w_500_223, w_500_224, w_500_225, w_500_226, w_500_227, w_500_228, w_500_229, w_500_230, w_500_231, w_500_232, w_500_233, w_500_234, w_500_235, w_500_236, w_500_237, w_500_238, w_500_239, w_500_240, w_500_241, w_500_242, w_500_243, w_500_244, w_500_245, w_500_246, w_500_247, w_500_248, w_500_249, w_500_250, w_500_251, w_500_252, w_500_253, w_500_254, w_500_255, w_500_256, w_500_257, w_500_258, w_500_259, w_500_260, w_500_261, w_500_262, w_500_263, w_500_264, w_500_265, w_500_266, w_500_267, w_500_268, w_500_269, w_500_270, w_500_271, w_500_272, w_500_273, w_500_274, w_500_275, w_500_276, w_500_277, w_500_278, w_500_279, w_500_280, w_500_281, w_500_282, w_500_283, w_500_284, w_500_285, w_500_286, w_500_287, w_500_288, w_500_289, w_500_290, w_500_291, w_500_292, w_500_293, w_500_294, w_500_295, w_500_296, w_500_297, w_500_298, w_500_299, w_500_300, w_500_301, w_500_302, w_500_303, w_500_304, w_500_305, w_500_306, w_500_307, w_500_308, w_500_309, w_500_310, w_500_311, w_500_312, w_500_313, w_500_314, w_500_315, w_500_316, w_500_317, w_500_318, w_500_319, w_500_320, w_500_321, w_500_322, w_500_323, w_500_324, w_500_325, w_500_326, w_500_327, w_500_328, w_500_329, w_500_330, w_500_331, w_500_332, w_500_333, w_500_334, w_500_335, w_500_336, w_500_337, w_500_338, w_500_339, w_500_340, w_500_341, w_500_342, w_500_343, w_500_344, w_500_345, w_500_346, w_500_347, w_500_348, w_500_349, w_500_350, w_500_351, w_500_352, w_500_353, w_500_354, w_500_355, w_500_356, w_500_357, w_500_358, w_500_359, w_500_360, w_500_361, w_500_362, w_500_363, w_500_364, w_500_365, w_500_366, w_500_367, w_500_368, w_500_369, w_500_370, w_500_371, w_500_372, w_500_373, w_500_374, w_500_375, w_500_376, w_500_377, w_500_378, w_500_379, w_500_380, w_500_381, w_500_382, w_500_383, w_500_384, w_500_385, w_500_386, w_500_387, w_500_388, w_500_389, w_500_390, w_500_391, w_500_392, w_500_393, w_500_394, w_500_395, w_500_396, w_500_397, w_500_398, w_500_399, w_500_400, w_500_401, w_500_402, w_500_403, w_500_404, w_500_405, w_500_406, w_500_407, w_500_408, w_500_409, w_500_410, w_500_411, w_500_412, w_500_413, w_500_414, w_500_415, w_500_416, w_500_417, w_500_418, w_500_419, w_500_420, w_500_421, w_500_422, w_500_423, w_500_424, w_500_425, w_500_426, w_500_427, w_500_428, w_500_429, w_500_430, w_500_431, w_500_432, w_500_433, w_500_434, w_500_435, w_500_436, w_500_437, w_500_438, w_500_439, w_500_440, w_500_441, w_500_442, w_500_443, w_500_444, w_500_445, w_500_446, w_500_447, w_500_448, w_500_449, w_500_450, w_500_451, w_500_452, w_500_453, w_500_454, w_500_455, w_500_456, w_500_457, w_500_458, w_500_459, w_500_460, w_500_461, w_500_462, w_500_463, w_500_464  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, r35, r36, r37, r38, r39, r40, r41, r42, r43, r44, r45, r46, r47, r48, r49, r50, r51, r52, r53, r54, r55, r56, r57, r58, r59, r60, r61, r62, r63, r64, r65, r66, r67, r68, r69, r70, r71, r72, r73, r74, r75, r76, r77, r78, r79, r80, r81, r82, r83, r84, r85, r86, r87, r88, r89, r90, r91, r92, r93, r94, r95, r96, r97, r98, r99, r100, r101, r102, r103, r104, r105, r106, r107, r108, r109, r110, r111, r112, r113, r114, r115, r116, r117, r118, r119, r120, r121, r122, r123, r124, r125, r126, r127, r128, r129, r130, r131, r132, r133, r134, r135, r136, r137, r138, r139, r140, r141, r142, r143, r144, r145, r146, r147, r148, r149, r150, r151, r152, r153, r154, r155, r156, r157, r158, r159, r160, r161, r162, r163, r164, r165, r166, r167, r168, r169, r170, r171, r172, r173, r174, r175, r176, r177, r178, r179, r180, r181, r182, r183, r184, r185, r186, r187, r188, r189, r190, r191, r192, r193, r194, r195, r196, r197, r198, r199, r200, r201, r202, r203, r204, r205, r206, r207, r208, r209, r210, r211, r212, r213, r214, r215, r216, r217, r218, r219, r220, r221, r222, r223, r224, r225, r226, r227, r228, r229, r230, r231, r232, r233, r234, r235, r236, r237, r238, r239, r240, r241, r242, r243, r244, r245, r246, r247, r248, r249, r250, r251, r252, r253, r254, r255, r256, r257, r258, r259, r260, r261, r262, r263, r264, r265, r266, r267, r268, r269, r270, r271, r272, r273, r274, r275, r276, r277, r278, r279, r280, r281, r282, r283, r284, r285, r286, r287, r288, r289, r290, r291, r292, r293, r294, r295, r296, r297, r298, r299, r300, r301, r302, r303, r304, r305, r306, r307, r308, r309, r310, r311, r312, r313, r314, r315, r316, r317, r318, r319, r320, r321, r322, r323, r324, r325, r326, r327, r328, r329, r330, r331, r332, r333, r334, r335, r336, r337, r338, r339, r340, r341, r342, r343, r344, r345, r346, r347, r348, r349, r350, r351, r352, r353, r354, r355, r356, r357, r358, r359, r360, r361, r362, r363, r364, r365, r366, r367, r368, r369, r370, r371, r372, r373, r374, r375, r376, r377, r378, r379, r380, r381, r382, r383, r384, r385, r386, r387, r388, r389, r390, r391, r392, r393, r394, r395, r396, r397, r398, r399, r400, r401, r402, r403, r404, r405, r406, r407, r408, r409, r410, r411, r412, r413, r414, r415, r416, r417, r418, r419, r420, r421, r422, r423, r424, r425, r426, r427, r428, r429, r430, r431, r432, r433, r434, r435, r436, r437, r438, r439, r440, r441, r442, r443, r444, r445, r446, r447, r448, r449, r450, r451, r452, r453, r454, r455, r456, r457, r458, r459, r460, r461, r462, r463, r464, r465, r466, r467, r468, r469, r470, r471, r472, r473, r474, r475, r476, r477, r478, r479, r480, r481, r482, r483, r484, r485, r486, r487, r488, r489, r490, r491, r492, r493, r494, r495, r496, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;
  assign w_000_035 = r35;
  assign w_000_036 = r36;
  assign w_000_037 = r37;
  assign w_000_038 = r38;
  assign w_000_039 = r39;
  assign w_000_040 = r40;
  assign w_000_041 = r41;
  assign w_000_042 = r42;
  assign w_000_043 = r43;
  assign w_000_044 = r44;
  assign w_000_045 = r45;
  assign w_000_046 = r46;
  assign w_000_047 = r47;
  assign w_000_048 = r48;
  assign w_000_049 = r49;
  assign w_000_050 = r50;
  assign w_000_051 = r51;
  assign w_000_052 = r52;
  assign w_000_053 = r53;
  assign w_000_054 = r54;
  assign w_000_055 = r55;
  assign w_000_056 = r56;
  assign w_000_057 = r57;
  assign w_000_058 = r58;
  assign w_000_059 = r59;
  assign w_000_060 = r60;
  assign w_000_061 = r61;
  assign w_000_062 = r62;
  assign w_000_063 = r63;
  assign w_000_064 = r64;
  assign w_000_065 = r65;
  assign w_000_066 = r66;
  assign w_000_067 = r67;
  assign w_000_068 = r68;
  assign w_000_069 = r69;
  assign w_000_070 = r70;
  assign w_000_071 = r71;
  assign w_000_072 = r72;
  assign w_000_073 = r73;
  assign w_000_074 = r74;
  assign w_000_075 = r75;
  assign w_000_076 = r76;
  assign w_000_077 = r77;
  assign w_000_078 = r78;
  assign w_000_079 = r79;
  assign w_000_080 = r80;
  assign w_000_081 = r81;
  assign w_000_082 = r82;
  assign w_000_083 = r83;
  assign w_000_084 = r84;
  assign w_000_085 = r85;
  assign w_000_086 = r86;
  assign w_000_087 = r87;
  assign w_000_088 = r88;
  assign w_000_089 = r89;
  assign w_000_090 = r90;
  assign w_000_091 = r91;
  assign w_000_092 = r92;
  assign w_000_093 = r93;
  assign w_000_094 = r94;
  assign w_000_095 = r95;
  assign w_000_096 = r96;
  assign w_000_097 = r97;
  assign w_000_098 = r98;
  assign w_000_099 = r99;
  assign w_000_100 = r100;
  assign w_000_101 = r101;
  assign w_000_102 = r102;
  assign w_000_103 = r103;
  assign w_000_104 = r104;
  assign w_000_105 = r105;
  assign w_000_106 = r106;
  assign w_000_107 = r107;
  assign w_000_108 = r108;
  assign w_000_109 = r109;
  assign w_000_110 = r110;
  assign w_000_111 = r111;
  assign w_000_112 = r112;
  assign w_000_113 = r113;
  assign w_000_114 = r114;
  assign w_000_115 = r115;
  assign w_000_116 = r116;
  assign w_000_117 = r117;
  assign w_000_118 = r118;
  assign w_000_119 = r119;
  assign w_000_120 = r120;
  assign w_000_121 = r121;
  assign w_000_122 = r122;
  assign w_000_123 = r123;
  assign w_000_124 = r124;
  assign w_000_125 = r125;
  assign w_000_126 = r126;
  assign w_000_127 = r127;
  assign w_000_128 = r128;
  assign w_000_129 = r129;
  assign w_000_130 = r130;
  assign w_000_131 = r131;
  assign w_000_132 = r132;
  assign w_000_133 = r133;
  assign w_000_134 = r134;
  assign w_000_135 = r135;
  assign w_000_136 = r136;
  assign w_000_137 = r137;
  assign w_000_138 = r138;
  assign w_000_139 = r139;
  assign w_000_140 = r140;
  assign w_000_141 = r141;
  assign w_000_142 = r142;
  assign w_000_143 = r143;
  assign w_000_144 = r144;
  assign w_000_145 = r145;
  assign w_000_146 = r146;
  assign w_000_147 = r147;
  assign w_000_148 = r148;
  assign w_000_149 = r149;
  assign w_000_150 = r150;
  assign w_000_151 = r151;
  assign w_000_152 = r152;
  assign w_000_153 = r153;
  assign w_000_154 = r154;
  assign w_000_155 = r155;
  assign w_000_156 = r156;
  assign w_000_157 = r157;
  assign w_000_158 = r158;
  assign w_000_159 = r159;
  assign w_000_160 = r160;
  assign w_000_161 = r161;
  assign w_000_162 = r162;
  assign w_000_163 = r163;
  assign w_000_164 = r164;
  assign w_000_165 = r165;
  assign w_000_166 = r166;
  assign w_000_167 = r167;
  assign w_000_168 = r168;
  assign w_000_169 = r169;
  assign w_000_170 = r170;
  assign w_000_171 = r171;
  assign w_000_172 = r172;
  assign w_000_173 = r173;
  assign w_000_174 = r174;
  assign w_000_175 = r175;
  assign w_000_176 = r176;
  assign w_000_177 = r177;
  assign w_000_178 = r178;
  assign w_000_179 = r179;
  assign w_000_180 = r180;
  assign w_000_181 = r181;
  assign w_000_182 = r182;
  assign w_000_183 = r183;
  assign w_000_184 = r184;
  assign w_000_185 = r185;
  assign w_000_186 = r186;
  assign w_000_187 = r187;
  assign w_000_188 = r188;
  assign w_000_189 = r189;
  assign w_000_190 = r190;
  assign w_000_191 = r191;
  assign w_000_192 = r192;
  assign w_000_193 = r193;
  assign w_000_194 = r194;
  assign w_000_195 = r195;
  assign w_000_196 = r196;
  assign w_000_197 = r197;
  assign w_000_198 = r198;
  assign w_000_199 = r199;
  assign w_000_200 = r200;
  assign w_000_201 = r201;
  assign w_000_202 = r202;
  assign w_000_203 = r203;
  assign w_000_204 = r204;
  assign w_000_205 = r205;
  assign w_000_206 = r206;
  assign w_000_207 = r207;
  assign w_000_208 = r208;
  assign w_000_209 = r209;
  assign w_000_210 = r210;
  assign w_000_211 = r211;
  assign w_000_212 = r212;
  assign w_000_213 = r213;
  assign w_000_214 = r214;
  assign w_000_215 = r215;
  assign w_000_216 = r216;
  assign w_000_217 = r217;
  assign w_000_218 = r218;
  assign w_000_219 = r219;
  assign w_000_220 = r220;
  assign w_000_221 = r221;
  assign w_000_222 = r222;
  assign w_000_223 = r223;
  assign w_000_224 = r224;
  assign w_000_225 = r225;
  assign w_000_226 = r226;
  assign w_000_227 = r227;
  assign w_000_228 = r228;
  assign w_000_229 = r229;
  assign w_000_230 = r230;
  assign w_000_231 = r231;
  assign w_000_232 = r232;
  assign w_000_233 = r233;
  assign w_000_234 = r234;
  assign w_000_235 = r235;
  assign w_000_236 = r236;
  assign w_000_237 = r237;
  assign w_000_238 = r238;
  assign w_000_239 = r239;
  assign w_000_240 = r240;
  assign w_000_241 = r241;
  assign w_000_242 = r242;
  assign w_000_243 = r243;
  assign w_000_244 = r244;
  assign w_000_245 = r245;
  assign w_000_246 = r246;
  assign w_000_247 = r247;
  assign w_000_248 = r248;
  assign w_000_249 = r249;
  assign w_000_250 = r250;
  assign w_000_251 = r251;
  assign w_000_252 = r252;
  assign w_000_253 = r253;
  assign w_000_254 = r254;
  assign w_000_255 = r255;
  assign w_000_256 = r256;
  assign w_000_257 = r257;
  assign w_000_258 = r258;
  assign w_000_259 = r259;
  assign w_000_260 = r260;
  assign w_000_261 = r261;
  assign w_000_262 = r262;
  assign w_000_263 = r263;
  assign w_000_264 = r264;
  assign w_000_265 = r265;
  assign w_000_266 = r266;
  assign w_000_267 = r267;
  assign w_000_268 = r268;
  assign w_000_269 = r269;
  assign w_000_270 = r270;
  assign w_000_271 = r271;
  assign w_000_272 = r272;
  assign w_000_273 = r273;
  assign w_000_274 = r274;
  assign w_000_275 = r275;
  assign w_000_276 = r276;
  assign w_000_277 = r277;
  assign w_000_278 = r278;
  assign w_000_279 = r279;
  assign w_000_280 = r280;
  assign w_000_281 = r281;
  assign w_000_282 = r282;
  assign w_000_283 = r283;
  assign w_000_284 = r284;
  assign w_000_285 = r285;
  assign w_000_286 = r286;
  assign w_000_287 = r287;
  assign w_000_288 = r288;
  assign w_000_289 = r289;
  assign w_000_290 = r290;
  assign w_000_291 = r291;
  assign w_000_292 = r292;
  assign w_000_293 = r293;
  assign w_000_294 = r294;
  assign w_000_295 = r295;
  assign w_000_296 = r296;
  assign w_000_297 = r297;
  assign w_000_298 = r298;
  assign w_000_299 = r299;
  assign w_000_300 = r300;
  assign w_000_301 = r301;
  assign w_000_302 = r302;
  assign w_000_303 = r303;
  assign w_000_304 = r304;
  assign w_000_305 = r305;
  assign w_000_306 = r306;
  assign w_000_307 = r307;
  assign w_000_308 = r308;
  assign w_000_309 = r309;
  assign w_000_310 = r310;
  assign w_000_311 = r311;
  assign w_000_312 = r312;
  assign w_000_313 = r313;
  assign w_000_314 = r314;
  assign w_000_315 = r315;
  assign w_000_316 = r316;
  assign w_000_317 = r317;
  assign w_000_318 = r318;
  assign w_000_319 = r319;
  assign w_000_320 = r320;
  assign w_000_321 = r321;
  assign w_000_322 = r322;
  assign w_000_323 = r323;
  assign w_000_324 = r324;
  assign w_000_325 = r325;
  assign w_000_326 = r326;
  assign w_000_327 = r327;
  assign w_000_328 = r328;
  assign w_000_329 = r329;
  assign w_000_330 = r330;
  assign w_000_331 = r331;
  assign w_000_332 = r332;
  assign w_000_333 = r333;
  assign w_000_334 = r334;
  assign w_000_335 = r335;
  assign w_000_336 = r336;
  assign w_000_337 = r337;
  assign w_000_338 = r338;
  assign w_000_339 = r339;
  assign w_000_340 = r340;
  assign w_000_341 = r341;
  assign w_000_342 = r342;
  assign w_000_343 = r343;
  assign w_000_344 = r344;
  assign w_000_345 = r345;
  assign w_000_346 = r346;
  assign w_000_347 = r347;
  assign w_000_348 = r348;
  assign w_000_349 = r349;
  assign w_000_350 = r350;
  assign w_000_351 = r351;
  assign w_000_352 = r352;
  assign w_000_353 = r353;
  assign w_000_354 = r354;
  assign w_000_355 = r355;
  assign w_000_356 = r356;
  assign w_000_357 = r357;
  assign w_000_358 = r358;
  assign w_000_359 = r359;
  assign w_000_360 = r360;
  assign w_000_361 = r361;
  assign w_000_362 = r362;
  assign w_000_363 = r363;
  assign w_000_364 = r364;
  assign w_000_365 = r365;
  assign w_000_366 = r366;
  assign w_000_367 = r367;
  assign w_000_368 = r368;
  assign w_000_369 = r369;
  assign w_000_370 = r370;
  assign w_000_371 = r371;
  assign w_000_372 = r372;
  assign w_000_373 = r373;
  assign w_000_374 = r374;
  assign w_000_375 = r375;
  assign w_000_376 = r376;
  assign w_000_377 = r377;
  assign w_000_378 = r378;
  assign w_000_379 = r379;
  assign w_000_380 = r380;
  assign w_000_381 = r381;
  assign w_000_382 = r382;
  assign w_000_383 = r383;
  assign w_000_384 = r384;
  assign w_000_385 = r385;
  assign w_000_386 = r386;
  assign w_000_387 = r387;
  assign w_000_388 = r388;
  assign w_000_389 = r389;
  assign w_000_390 = r390;
  assign w_000_391 = r391;
  assign w_000_392 = r392;
  assign w_000_393 = r393;
  assign w_000_394 = r394;
  assign w_000_395 = r395;
  assign w_000_396 = r396;
  assign w_000_397 = r397;
  assign w_000_398 = r398;
  assign w_000_399 = r399;
  assign w_000_400 = r400;
  assign w_000_401 = r401;
  assign w_000_402 = r402;
  assign w_000_403 = r403;
  assign w_000_404 = r404;
  assign w_000_405 = r405;
  assign w_000_406 = r406;
  assign w_000_407 = r407;
  assign w_000_408 = r408;
  assign w_000_409 = r409;
  assign w_000_410 = r410;
  assign w_000_411 = r411;
  assign w_000_412 = r412;
  assign w_000_413 = r413;
  assign w_000_414 = r414;
  assign w_000_415 = r415;
  assign w_000_416 = r416;
  assign w_000_417 = r417;
  assign w_000_418 = r418;
  assign w_000_419 = r419;
  assign w_000_420 = r420;
  assign w_000_421 = r421;
  assign w_000_422 = r422;
  assign w_000_423 = r423;
  assign w_000_424 = r424;
  assign w_000_425 = r425;
  assign w_000_426 = r426;
  assign w_000_427 = r427;
  assign w_000_428 = r428;
  assign w_000_429 = r429;
  assign w_000_430 = r430;
  assign w_000_431 = r431;
  assign w_000_432 = r432;
  assign w_000_433 = r433;
  assign w_000_434 = r434;
  assign w_000_435 = r435;
  assign w_000_436 = r436;
  assign w_000_437 = r437;
  assign w_000_438 = r438;
  assign w_000_439 = r439;
  assign w_000_440 = r440;
  assign w_000_441 = r441;
  assign w_000_442 = r442;
  assign w_000_443 = r443;
  assign w_000_444 = r444;
  assign w_000_445 = r445;
  assign w_000_446 = r446;
  assign w_000_447 = r447;
  assign w_000_448 = r448;
  assign w_000_449 = r449;
  assign w_000_450 = r450;
  assign w_000_451 = r451;
  assign w_000_452 = r452;
  assign w_000_453 = r453;
  assign w_000_454 = r454;
  assign w_000_455 = r455;
  assign w_000_456 = r456;
  assign w_000_457 = r457;
  assign w_000_458 = r458;
  assign w_000_459 = r459;
  assign w_000_460 = r460;
  assign w_000_461 = r461;
  assign w_000_462 = r462;
  assign w_000_463 = r463;
  assign w_000_464 = r464;
  assign w_000_465 = r465;
  assign w_000_466 = r466;
  assign w_000_467 = r467;
  assign w_000_468 = r468;
  assign w_000_469 = r469;
  assign w_000_470 = r470;
  assign w_000_471 = r471;
  assign w_000_472 = r472;
  assign w_000_473 = r473;
  assign w_000_474 = r474;
  assign w_000_475 = r475;
  assign w_000_476 = r476;
  assign w_000_477 = r477;
  assign w_000_478 = r478;
  assign w_000_479 = r479;
  assign w_000_480 = r480;
  assign w_000_481 = r481;
  assign w_000_482 = r482;
  assign w_000_483 = r483;
  assign w_000_484 = r484;
  assign w_000_485 = r485;
  assign w_000_486 = r486;
  assign w_000_487 = r487;
  assign w_000_488 = r488;
  assign w_000_489 = r489;
  assign w_000_490 = r490;
  assign w_000_491 = r491;
  assign w_000_492 = r492;
  assign w_000_493 = r493;
  assign w_000_494 = r494;
  assign w_000_495 = r495;
  assign w_000_496 = r496;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    r35 = 1'b0; 
    r36 = 1'b0; 
    r37 = 1'b0; 
    r38 = 1'b0; 
    r39 = 1'b0; 
    r40 = 1'b0; 
    r41 = 1'b0; 
    r42 = 1'b0; 
    r43 = 1'b0; 
    r44 = 1'b0; 
    r45 = 1'b0; 
    r46 = 1'b0; 
    r47 = 1'b0; 
    r48 = 1'b0; 
    r49 = 1'b0; 
    r50 = 1'b0; 
    r51 = 1'b0; 
    r52 = 1'b0; 
    r53 = 1'b0; 
    r54 = 1'b0; 
    r55 = 1'b0; 
    r56 = 1'b0; 
    r57 = 1'b0; 
    r58 = 1'b0; 
    r59 = 1'b0; 
    r60 = 1'b0; 
    r61 = 1'b0; 
    r62 = 1'b0; 
    r63 = 1'b0; 
    r64 = 1'b0; 
    r65 = 1'b0; 
    r66 = 1'b0; 
    r67 = 1'b0; 
    r68 = 1'b0; 
    r69 = 1'b0; 
    r70 = 1'b0; 
    r71 = 1'b0; 
    r72 = 1'b0; 
    r73 = 1'b0; 
    r74 = 1'b0; 
    r75 = 1'b0; 
    r76 = 1'b0; 
    r77 = 1'b0; 
    r78 = 1'b0; 
    r79 = 1'b0; 
    r80 = 1'b0; 
    r81 = 1'b0; 
    r82 = 1'b0; 
    r83 = 1'b0; 
    r84 = 1'b0; 
    r85 = 1'b0; 
    r86 = 1'b0; 
    r87 = 1'b0; 
    r88 = 1'b0; 
    r89 = 1'b0; 
    r90 = 1'b0; 
    r91 = 1'b0; 
    r92 = 1'b0; 
    r93 = 1'b0; 
    r94 = 1'b0; 
    r95 = 1'b0; 
    r96 = 1'b0; 
    r97 = 1'b0; 
    r98 = 1'b0; 
    r99 = 1'b0; 
    r100 = 1'b0; 
    r101 = 1'b0; 
    r102 = 1'b0; 
    r103 = 1'b0; 
    r104 = 1'b0; 
    r105 = 1'b0; 
    r106 = 1'b0; 
    r107 = 1'b0; 
    r108 = 1'b0; 
    r109 = 1'b0; 
    r110 = 1'b0; 
    r111 = 1'b0; 
    r112 = 1'b0; 
    r113 = 1'b0; 
    r114 = 1'b0; 
    r115 = 1'b0; 
    r116 = 1'b0; 
    r117 = 1'b0; 
    r118 = 1'b0; 
    r119 = 1'b0; 
    r120 = 1'b0; 
    r121 = 1'b0; 
    r122 = 1'b0; 
    r123 = 1'b0; 
    r124 = 1'b0; 
    r125 = 1'b0; 
    r126 = 1'b0; 
    r127 = 1'b0; 
    r128 = 1'b0; 
    r129 = 1'b0; 
    r130 = 1'b0; 
    r131 = 1'b0; 
    r132 = 1'b0; 
    r133 = 1'b0; 
    r134 = 1'b0; 
    r135 = 1'b0; 
    r136 = 1'b0; 
    r137 = 1'b0; 
    r138 = 1'b0; 
    r139 = 1'b0; 
    r140 = 1'b0; 
    r141 = 1'b0; 
    r142 = 1'b0; 
    r143 = 1'b0; 
    r144 = 1'b0; 
    r145 = 1'b0; 
    r146 = 1'b0; 
    r147 = 1'b0; 
    r148 = 1'b0; 
    r149 = 1'b0; 
    r150 = 1'b0; 
    r151 = 1'b0; 
    r152 = 1'b0; 
    r153 = 1'b0; 
    r154 = 1'b0; 
    r155 = 1'b0; 
    r156 = 1'b0; 
    r157 = 1'b0; 
    r158 = 1'b0; 
    r159 = 1'b0; 
    r160 = 1'b0; 
    r161 = 1'b0; 
    r162 = 1'b0; 
    r163 = 1'b0; 
    r164 = 1'b0; 
    r165 = 1'b0; 
    r166 = 1'b0; 
    r167 = 1'b0; 
    r168 = 1'b0; 
    r169 = 1'b0; 
    r170 = 1'b0; 
    r171 = 1'b0; 
    r172 = 1'b0; 
    r173 = 1'b0; 
    r174 = 1'b0; 
    r175 = 1'b0; 
    r176 = 1'b0; 
    r177 = 1'b0; 
    r178 = 1'b0; 
    r179 = 1'b0; 
    r180 = 1'b0; 
    r181 = 1'b0; 
    r182 = 1'b0; 
    r183 = 1'b0; 
    r184 = 1'b0; 
    r185 = 1'b0; 
    r186 = 1'b0; 
    r187 = 1'b0; 
    r188 = 1'b0; 
    r189 = 1'b0; 
    r190 = 1'b0; 
    r191 = 1'b0; 
    r192 = 1'b0; 
    r193 = 1'b0; 
    r194 = 1'b0; 
    r195 = 1'b0; 
    r196 = 1'b0; 
    r197 = 1'b0; 
    r198 = 1'b0; 
    r199 = 1'b0; 
    r200 = 1'b0; 
    r201 = 1'b0; 
    r202 = 1'b0; 
    r203 = 1'b0; 
    r204 = 1'b0; 
    r205 = 1'b0; 
    r206 = 1'b0; 
    r207 = 1'b0; 
    r208 = 1'b0; 
    r209 = 1'b0; 
    r210 = 1'b0; 
    r211 = 1'b0; 
    r212 = 1'b0; 
    r213 = 1'b0; 
    r214 = 1'b0; 
    r215 = 1'b0; 
    r216 = 1'b0; 
    r217 = 1'b0; 
    r218 = 1'b0; 
    r219 = 1'b0; 
    r220 = 1'b0; 
    r221 = 1'b0; 
    r222 = 1'b0; 
    r223 = 1'b0; 
    r224 = 1'b0; 
    r225 = 1'b0; 
    r226 = 1'b0; 
    r227 = 1'b0; 
    r228 = 1'b0; 
    r229 = 1'b0; 
    r230 = 1'b0; 
    r231 = 1'b0; 
    r232 = 1'b0; 
    r233 = 1'b0; 
    r234 = 1'b0; 
    r235 = 1'b0; 
    r236 = 1'b0; 
    r237 = 1'b0; 
    r238 = 1'b0; 
    r239 = 1'b0; 
    r240 = 1'b0; 
    r241 = 1'b0; 
    r242 = 1'b0; 
    r243 = 1'b0; 
    r244 = 1'b0; 
    r245 = 1'b0; 
    r246 = 1'b0; 
    r247 = 1'b0; 
    r248 = 1'b0; 
    r249 = 1'b0; 
    r250 = 1'b0; 
    r251 = 1'b0; 
    r252 = 1'b0; 
    r253 = 1'b0; 
    r254 = 1'b0; 
    r255 = 1'b0; 
    r256 = 1'b0; 
    r257 = 1'b0; 
    r258 = 1'b0; 
    r259 = 1'b0; 
    r260 = 1'b0; 
    r261 = 1'b0; 
    r262 = 1'b0; 
    r263 = 1'b0; 
    r264 = 1'b0; 
    r265 = 1'b0; 
    r266 = 1'b0; 
    r267 = 1'b0; 
    r268 = 1'b0; 
    r269 = 1'b0; 
    r270 = 1'b0; 
    r271 = 1'b0; 
    r272 = 1'b0; 
    r273 = 1'b0; 
    r274 = 1'b0; 
    r275 = 1'b0; 
    r276 = 1'b0; 
    r277 = 1'b0; 
    r278 = 1'b0; 
    r279 = 1'b0; 
    r280 = 1'b0; 
    r281 = 1'b0; 
    r282 = 1'b0; 
    r283 = 1'b0; 
    r284 = 1'b0; 
    r285 = 1'b0; 
    r286 = 1'b0; 
    r287 = 1'b0; 
    r288 = 1'b0; 
    r289 = 1'b0; 
    r290 = 1'b0; 
    r291 = 1'b0; 
    r292 = 1'b0; 
    r293 = 1'b0; 
    r294 = 1'b0; 
    r295 = 1'b0; 
    r296 = 1'b0; 
    r297 = 1'b0; 
    r298 = 1'b0; 
    r299 = 1'b0; 
    r300 = 1'b0; 
    r301 = 1'b0; 
    r302 = 1'b0; 
    r303 = 1'b0; 
    r304 = 1'b0; 
    r305 = 1'b0; 
    r306 = 1'b0; 
    r307 = 1'b0; 
    r308 = 1'b0; 
    r309 = 1'b0; 
    r310 = 1'b0; 
    r311 = 1'b0; 
    r312 = 1'b0; 
    r313 = 1'b0; 
    r314 = 1'b0; 
    r315 = 1'b0; 
    r316 = 1'b0; 
    r317 = 1'b0; 
    r318 = 1'b0; 
    r319 = 1'b0; 
    r320 = 1'b0; 
    r321 = 1'b0; 
    r322 = 1'b0; 
    r323 = 1'b0; 
    r324 = 1'b0; 
    r325 = 1'b0; 
    r326 = 1'b0; 
    r327 = 1'b0; 
    r328 = 1'b0; 
    r329 = 1'b0; 
    r330 = 1'b0; 
    r331 = 1'b0; 
    r332 = 1'b0; 
    r333 = 1'b0; 
    r334 = 1'b0; 
    r335 = 1'b0; 
    r336 = 1'b0; 
    r337 = 1'b0; 
    r338 = 1'b0; 
    r339 = 1'b0; 
    r340 = 1'b0; 
    r341 = 1'b0; 
    r342 = 1'b0; 
    r343 = 1'b0; 
    r344 = 1'b0; 
    r345 = 1'b0; 
    r346 = 1'b0; 
    r347 = 1'b0; 
    r348 = 1'b0; 
    r349 = 1'b0; 
    r350 = 1'b0; 
    r351 = 1'b0; 
    r352 = 1'b0; 
    r353 = 1'b0; 
    r354 = 1'b0; 
    r355 = 1'b0; 
    r356 = 1'b0; 
    r357 = 1'b0; 
    r358 = 1'b0; 
    r359 = 1'b0; 
    r360 = 1'b0; 
    r361 = 1'b0; 
    r362 = 1'b0; 
    r363 = 1'b0; 
    r364 = 1'b0; 
    r365 = 1'b0; 
    r366 = 1'b0; 
    r367 = 1'b0; 
    r368 = 1'b0; 
    r369 = 1'b0; 
    r370 = 1'b0; 
    r371 = 1'b0; 
    r372 = 1'b0; 
    r373 = 1'b0; 
    r374 = 1'b0; 
    r375 = 1'b0; 
    r376 = 1'b0; 
    r377 = 1'b0; 
    r378 = 1'b0; 
    r379 = 1'b0; 
    r380 = 1'b0; 
    r381 = 1'b0; 
    r382 = 1'b0; 
    r383 = 1'b0; 
    r384 = 1'b0; 
    r385 = 1'b0; 
    r386 = 1'b0; 
    r387 = 1'b0; 
    r388 = 1'b0; 
    r389 = 1'b0; 
    r390 = 1'b0; 
    r391 = 1'b0; 
    r392 = 1'b0; 
    r393 = 1'b0; 
    r394 = 1'b0; 
    r395 = 1'b0; 
    r396 = 1'b0; 
    r397 = 1'b0; 
    r398 = 1'b0; 
    r399 = 1'b0; 
    r400 = 1'b0; 
    r401 = 1'b0; 
    r402 = 1'b0; 
    r403 = 1'b0; 
    r404 = 1'b0; 
    r405 = 1'b0; 
    r406 = 1'b0; 
    r407 = 1'b0; 
    r408 = 1'b0; 
    r409 = 1'b0; 
    r410 = 1'b0; 
    r411 = 1'b0; 
    r412 = 1'b0; 
    r413 = 1'b0; 
    r414 = 1'b0; 
    r415 = 1'b0; 
    r416 = 1'b0; 
    r417 = 1'b0; 
    r418 = 1'b0; 
    r419 = 1'b0; 
    r420 = 1'b0; 
    r421 = 1'b0; 
    r422 = 1'b0; 
    r423 = 1'b0; 
    r424 = 1'b0; 
    r425 = 1'b0; 
    r426 = 1'b0; 
    r427 = 1'b0; 
    r428 = 1'b0; 
    r429 = 1'b0; 
    r430 = 1'b0; 
    r431 = 1'b0; 
    r432 = 1'b0; 
    r433 = 1'b0; 
    r434 = 1'b0; 
    r435 = 1'b0; 
    r436 = 1'b0; 
    r437 = 1'b0; 
    r438 = 1'b0; 
    r439 = 1'b0; 
    r440 = 1'b0; 
    r441 = 1'b0; 
    r442 = 1'b0; 
    r443 = 1'b0; 
    r444 = 1'b0; 
    r445 = 1'b0; 
    r446 = 1'b0; 
    r447 = 1'b0; 
    r448 = 1'b0; 
    r449 = 1'b0; 
    r450 = 1'b0; 
    r451 = 1'b0; 
    r452 = 1'b0; 
    r453 = 1'b0; 
    r454 = 1'b0; 
    r455 = 1'b0; 
    r456 = 1'b0; 
    r457 = 1'b0; 
    r458 = 1'b0; 
    r459 = 1'b0; 
    r460 = 1'b0; 
    r461 = 1'b0; 
    r462 = 1'b0; 
    r463 = 1'b0; 
    r464 = 1'b0; 
    r465 = 1'b0; 
    r466 = 1'b0; 
    r467 = 1'b0; 
    r468 = 1'b0; 
    r469 = 1'b0; 
    r470 = 1'b0; 
    r471 = 1'b0; 
    r472 = 1'b0; 
    r473 = 1'b0; 
    r474 = 1'b0; 
    r475 = 1'b0; 
    r476 = 1'b0; 
    r477 = 1'b0; 
    r478 = 1'b0; 
    r479 = 1'b0; 
    r480 = 1'b0; 
    r481 = 1'b0; 
    r482 = 1'b0; 
    r483 = 1'b0; 
    r484 = 1'b0; 
    r485 = 1'b0; 
    r486 = 1'b0; 
    r487 = 1'b0; 
    r488 = 1'b0; 
    r489 = 1'b0; 
    r490 = 1'b0; 
    r491 = 1'b0; 
    r492 = 1'b0; 
    r493 = 1'b0; 
    r494 = 1'b0; 
    r495 = 1'b0; 
    r496 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_500_000, w_500_001, w_500_002, w_500_003, w_500_004, w_500_005, w_500_006, w_500_007, w_500_008, w_500_009, w_500_010, w_500_011, w_500_012, w_500_013, w_500_014, w_500_015, w_500_016, w_500_017, w_500_018, w_500_019, w_500_020, w_500_021, w_500_022, w_500_023, w_500_024, w_500_025, w_500_026, w_500_027, w_500_028, w_500_029, w_500_030, w_500_031, w_500_032, w_500_033, w_500_034, w_500_035, w_500_036, w_500_037, w_500_038, w_500_039, w_500_040, w_500_041, w_500_042, w_500_043, w_500_044, w_500_045, w_500_046, w_500_047, w_500_048, w_500_049, w_500_050, w_500_051, w_500_052, w_500_053, w_500_054, w_500_055, w_500_056, w_500_057, w_500_058, w_500_059, w_500_060, w_500_061, w_500_062, w_500_063, w_500_064, w_500_065, w_500_066, w_500_067, w_500_068, w_500_069, w_500_070, w_500_071, w_500_072, w_500_073, w_500_074, w_500_075, w_500_076, w_500_077, w_500_078, w_500_079, w_500_080, w_500_081, w_500_082, w_500_083, w_500_084, w_500_085, w_500_086, w_500_087, w_500_088, w_500_089, w_500_090, w_500_091, w_500_092, w_500_093, w_500_094, w_500_095, w_500_096, w_500_097, w_500_098, w_500_099, w_500_100, w_500_101, w_500_102, w_500_103, w_500_104, w_500_105, w_500_106, w_500_107, w_500_108, w_500_109, w_500_110, w_500_111, w_500_112, w_500_113, w_500_114, w_500_115, w_500_116, w_500_117, w_500_118, w_500_119, w_500_120, w_500_121, w_500_122, w_500_123, w_500_124, w_500_125, w_500_126, w_500_127, w_500_128, w_500_129, w_500_130, w_500_131, w_500_132, w_500_133, w_500_134, w_500_135, w_500_136, w_500_137, w_500_138, w_500_139, w_500_140, w_500_141, w_500_142, w_500_143, w_500_144, w_500_145, w_500_146, w_500_147, w_500_148, w_500_149, w_500_150, w_500_151, w_500_152, w_500_153, w_500_154, w_500_155, w_500_156, w_500_157, w_500_158, w_500_159, w_500_160, w_500_161, w_500_162, w_500_163, w_500_164, w_500_165, w_500_166, w_500_167, w_500_168, w_500_169, w_500_170, w_500_171, w_500_172, w_500_173, w_500_174, w_500_175, w_500_176, w_500_177, w_500_178, w_500_179, w_500_180, w_500_181, w_500_182, w_500_183, w_500_184, w_500_185, w_500_186, w_500_187, w_500_188, w_500_189, w_500_190, w_500_191, w_500_192, w_500_193, w_500_194, w_500_195, w_500_196, w_500_197, w_500_198, w_500_199, w_500_200, w_500_201, w_500_202, w_500_203, w_500_204, w_500_205, w_500_206, w_500_207, w_500_208, w_500_209, w_500_210, w_500_211, w_500_212, w_500_213, w_500_214, w_500_215, w_500_216, w_500_217, w_500_218, w_500_219, w_500_220, w_500_221, w_500_222, w_500_223, w_500_224, w_500_225, w_500_226, w_500_227, w_500_228, w_500_229, w_500_230, w_500_231, w_500_232, w_500_233, w_500_234, w_500_235, w_500_236, w_500_237, w_500_238, w_500_239, w_500_240, w_500_241, w_500_242, w_500_243, w_500_244, w_500_245, w_500_246, w_500_247, w_500_248, w_500_249, w_500_250, w_500_251, w_500_252, w_500_253, w_500_254, w_500_255, w_500_256, w_500_257, w_500_258, w_500_259, w_500_260, w_500_261, w_500_262, w_500_263, w_500_264, w_500_265, w_500_266, w_500_267, w_500_268, w_500_269, w_500_270, w_500_271, w_500_272, w_500_273, w_500_274, w_500_275, w_500_276, w_500_277, w_500_278, w_500_279, w_500_280, w_500_281, w_500_282, w_500_283, w_500_284, w_500_285, w_500_286, w_500_287, w_500_288, w_500_289, w_500_290, w_500_291, w_500_292, w_500_293, w_500_294, w_500_295, w_500_296, w_500_297, w_500_298, w_500_299, w_500_300, w_500_301, w_500_302, w_500_303, w_500_304, w_500_305, w_500_306, w_500_307, w_500_308, w_500_309, w_500_310, w_500_311, w_500_312, w_500_313, w_500_314, w_500_315, w_500_316, w_500_317, w_500_318, w_500_319, w_500_320, w_500_321, w_500_322, w_500_323, w_500_324, w_500_325, w_500_326, w_500_327, w_500_328, w_500_329, w_500_330, w_500_331, w_500_332, w_500_333, w_500_334, w_500_335, w_500_336, w_500_337, w_500_338, w_500_339, w_500_340, w_500_341, w_500_342, w_500_343, w_500_344, w_500_345, w_500_346, w_500_347, w_500_348, w_500_349, w_500_350, w_500_351, w_500_352, w_500_353, w_500_354, w_500_355, w_500_356, w_500_357, w_500_358, w_500_359, w_500_360, w_500_361, w_500_362, w_500_363, w_500_364, w_500_365, w_500_366, w_500_367, w_500_368, w_500_369, w_500_370, w_500_371, w_500_372, w_500_373, w_500_374, w_500_375, w_500_376, w_500_377, w_500_378, w_500_379, w_500_380, w_500_381, w_500_382, w_500_383, w_500_384, w_500_385, w_500_386, w_500_387, w_500_388, w_500_389, w_500_390, w_500_391, w_500_392, w_500_393, w_500_394, w_500_395, w_500_396, w_500_397, w_500_398, w_500_399, w_500_400, w_500_401, w_500_402, w_500_403, w_500_404, w_500_405, w_500_406, w_500_407, w_500_408, w_500_409, w_500_410, w_500_411, w_500_412, w_500_413, w_500_414, w_500_415, w_500_416, w_500_417, w_500_418, w_500_419, w_500_420, w_500_421, w_500_422, w_500_423, w_500_424, w_500_425, w_500_426, w_500_427, w_500_428, w_500_429, w_500_430, w_500_431, w_500_432, w_500_433, w_500_434, w_500_435, w_500_436, w_500_437, w_500_438, w_500_439, w_500_440, w_500_441, w_500_442, w_500_443, w_500_444, w_500_445, w_500_446, w_500_447, w_500_448, w_500_449, w_500_450, w_500_451, w_500_452, w_500_453, w_500_454, w_500_455, w_500_456, w_500_457, w_500_458, w_500_459, w_500_460, w_500_461, w_500_462, w_500_463, w_500_464);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
  always #34359738368 r35 = ~r35;
  always #68719476736 r36 = ~r36;
  always #137438953472 r37 = ~r37;
  always #274877906944 r38 = ~r38;
  always #549755813888 r39 = ~r39;
  always #1099511627776 r40 = ~r40;
  always #2199023255552 r41 = ~r41;
  always #4398046511104 r42 = ~r42;
  always #8796093022208 r43 = ~r43;
  always #17592186044416 r44 = ~r44;
  always #35184372088832 r45 = ~r45;
  always #70368744177664 r46 = ~r46;
  always #140737488355328 r47 = ~r47;
  always #281474976710656 r48 = ~r48;
  always #562949953421312 r49 = ~r49;
  always #1125899906842624 r50 = ~r50;
  always #2251799813685248 r51 = ~r51;
  always #4503599627370496 r52 = ~r52;
  always #9007199254740992 r53 = ~r53;
  always #18014398509481984 r54 = ~r54;
  always #36028797018963968 r55 = ~r55;
  always #72057594037927936 r56 = ~r56;
  always #144115188075855872 r57 = ~r57;
  always #288230376151711744 r58 = ~r58;
  always #576460752303423488 r59 = ~r59;
  always #1152921504606846976 r60 = ~r60;
  always #2305843009213693952 r61 = ~r61;
  always #4611686018427387904 r62 = ~r62;
  always #9223372036854775808 r63 = ~r63;
  always #1 r64 = ~r64;
  always #2 r65 = ~r65;
  always #4 r66 = ~r66;
  always #8 r67 = ~r67;
  always #16 r68 = ~r68;
  always #32 r69 = ~r69;
  always #64 r70 = ~r70;
  always #128 r71 = ~r71;
  always #256 r72 = ~r72;
  always #512 r73 = ~r73;
  always #1024 r74 = ~r74;
  always #2048 r75 = ~r75;
  always #4096 r76 = ~r76;
  always #8192 r77 = ~r77;
  always #16384 r78 = ~r78;
  always #32768 r79 = ~r79;
  always #65536 r80 = ~r80;
  always #131072 r81 = ~r81;
  always #262144 r82 = ~r82;
  always #524288 r83 = ~r83;
  always #1048576 r84 = ~r84;
  always #2097152 r85 = ~r85;
  always #4194304 r86 = ~r86;
  always #8388608 r87 = ~r87;
  always #16777216 r88 = ~r88;
  always #33554432 r89 = ~r89;
  always #67108864 r90 = ~r90;
  always #134217728 r91 = ~r91;
  always #268435456 r92 = ~r92;
  always #536870912 r93 = ~r93;
  always #1073741824 r94 = ~r94;
  always #2147483648 r95 = ~r95;
  always #4294967296 r96 = ~r96;
  always #8589934592 r97 = ~r97;
  always #17179869184 r98 = ~r98;
  always #34359738368 r99 = ~r99;
  always #68719476736 r100 = ~r100;
  always #137438953472 r101 = ~r101;
  always #274877906944 r102 = ~r102;
  always #549755813888 r103 = ~r103;
  always #1099511627776 r104 = ~r104;
  always #2199023255552 r105 = ~r105;
  always #4398046511104 r106 = ~r106;
  always #8796093022208 r107 = ~r107;
  always #17592186044416 r108 = ~r108;
  always #35184372088832 r109 = ~r109;
  always #70368744177664 r110 = ~r110;
  always #140737488355328 r111 = ~r111;
  always #281474976710656 r112 = ~r112;
  always #562949953421312 r113 = ~r113;
  always #1125899906842624 r114 = ~r114;
  always #2251799813685248 r115 = ~r115;
  always #4503599627370496 r116 = ~r116;
  always #9007199254740992 r117 = ~r117;
  always #18014398509481984 r118 = ~r118;
  always #36028797018963968 r119 = ~r119;
  always #72057594037927936 r120 = ~r120;
  always #144115188075855872 r121 = ~r121;
  always #288230376151711744 r122 = ~r122;
  always #576460752303423488 r123 = ~r123;
  always #1152921504606846976 r124 = ~r124;
  always #2305843009213693952 r125 = ~r125;
  always #4611686018427387904 r126 = ~r126;
  always #9223372036854775808 r127 = ~r127;
  always #1 r128 = ~r128;
  always #2 r129 = ~r129;
  always #4 r130 = ~r130;
  always #8 r131 = ~r131;
  always #16 r132 = ~r132;
  always #32 r133 = ~r133;
  always #64 r134 = ~r134;
  always #128 r135 = ~r135;
  always #256 r136 = ~r136;
  always #512 r137 = ~r137;
  always #1024 r138 = ~r138;
  always #2048 r139 = ~r139;
  always #4096 r140 = ~r140;
  always #8192 r141 = ~r141;
  always #16384 r142 = ~r142;
  always #32768 r143 = ~r143;
  always #65536 r144 = ~r144;
  always #131072 r145 = ~r145;
  always #262144 r146 = ~r146;
  always #524288 r147 = ~r147;
  always #1048576 r148 = ~r148;
  always #2097152 r149 = ~r149;
  always #4194304 r150 = ~r150;
  always #8388608 r151 = ~r151;
  always #16777216 r152 = ~r152;
  always #33554432 r153 = ~r153;
  always #67108864 r154 = ~r154;
  always #134217728 r155 = ~r155;
  always #268435456 r156 = ~r156;
  always #536870912 r157 = ~r157;
  always #1073741824 r158 = ~r158;
  always #2147483648 r159 = ~r159;
  always #4294967296 r160 = ~r160;
  always #8589934592 r161 = ~r161;
  always #17179869184 r162 = ~r162;
  always #34359738368 r163 = ~r163;
  always #68719476736 r164 = ~r164;
  always #137438953472 r165 = ~r165;
  always #274877906944 r166 = ~r166;
  always #549755813888 r167 = ~r167;
  always #1099511627776 r168 = ~r168;
  always #2199023255552 r169 = ~r169;
  always #4398046511104 r170 = ~r170;
  always #8796093022208 r171 = ~r171;
  always #17592186044416 r172 = ~r172;
  always #35184372088832 r173 = ~r173;
  always #70368744177664 r174 = ~r174;
  always #140737488355328 r175 = ~r175;
  always #281474976710656 r176 = ~r176;
  always #562949953421312 r177 = ~r177;
  always #1125899906842624 r178 = ~r178;
  always #2251799813685248 r179 = ~r179;
  always #4503599627370496 r180 = ~r180;
  always #9007199254740992 r181 = ~r181;
  always #18014398509481984 r182 = ~r182;
  always #36028797018963968 r183 = ~r183;
  always #72057594037927936 r184 = ~r184;
  always #144115188075855872 r185 = ~r185;
  always #288230376151711744 r186 = ~r186;
  always #576460752303423488 r187 = ~r187;
  always #1152921504606846976 r188 = ~r188;
  always #2305843009213693952 r189 = ~r189;
  always #4611686018427387904 r190 = ~r190;
  always #9223372036854775808 r191 = ~r191;
  always #1 r192 = ~r192;
  always #2 r193 = ~r193;
  always #4 r194 = ~r194;
  always #8 r195 = ~r195;
  always #16 r196 = ~r196;
  always #32 r197 = ~r197;
  always #64 r198 = ~r198;
  always #128 r199 = ~r199;
  always #256 r200 = ~r200;
  always #512 r201 = ~r201;
  always #1024 r202 = ~r202;
  always #2048 r203 = ~r203;
  always #4096 r204 = ~r204;
  always #8192 r205 = ~r205;
  always #16384 r206 = ~r206;
  always #32768 r207 = ~r207;
  always #65536 r208 = ~r208;
  always #131072 r209 = ~r209;
  always #262144 r210 = ~r210;
  always #524288 r211 = ~r211;
  always #1048576 r212 = ~r212;
  always #2097152 r213 = ~r213;
  always #4194304 r214 = ~r214;
  always #8388608 r215 = ~r215;
  always #16777216 r216 = ~r216;
  always #33554432 r217 = ~r217;
  always #67108864 r218 = ~r218;
  always #134217728 r219 = ~r219;
  always #268435456 r220 = ~r220;
  always #536870912 r221 = ~r221;
  always #1073741824 r222 = ~r222;
  always #2147483648 r223 = ~r223;
  always #4294967296 r224 = ~r224;
  always #8589934592 r225 = ~r225;
  always #17179869184 r226 = ~r226;
  always #34359738368 r227 = ~r227;
  always #68719476736 r228 = ~r228;
  always #137438953472 r229 = ~r229;
  always #274877906944 r230 = ~r230;
  always #549755813888 r231 = ~r231;
  always #1099511627776 r232 = ~r232;
  always #2199023255552 r233 = ~r233;
  always #4398046511104 r234 = ~r234;
  always #8796093022208 r235 = ~r235;
  always #17592186044416 r236 = ~r236;
  always #35184372088832 r237 = ~r237;
  always #70368744177664 r238 = ~r238;
  always #140737488355328 r239 = ~r239;
  always #281474976710656 r240 = ~r240;
  always #562949953421312 r241 = ~r241;
  always #1125899906842624 r242 = ~r242;
  always #2251799813685248 r243 = ~r243;
  always #4503599627370496 r244 = ~r244;
  always #9007199254740992 r245 = ~r245;
  always #18014398509481984 r246 = ~r246;
  always #36028797018963968 r247 = ~r247;
  always #72057594037927936 r248 = ~r248;
  always #144115188075855872 r249 = ~r249;
  always #288230376151711744 r250 = ~r250;
  always #576460752303423488 r251 = ~r251;
  always #1152921504606846976 r252 = ~r252;
  always #2305843009213693952 r253 = ~r253;
  always #4611686018427387904 r254 = ~r254;
  always #9223372036854775808 r255 = ~r255;
  always #1 r256 = ~r256;
  always #2 r257 = ~r257;
  always #4 r258 = ~r258;
  always #8 r259 = ~r259;
  always #16 r260 = ~r260;
  always #32 r261 = ~r261;
  always #64 r262 = ~r262;
  always #128 r263 = ~r263;
  always #256 r264 = ~r264;
  always #512 r265 = ~r265;
  always #1024 r266 = ~r266;
  always #2048 r267 = ~r267;
  always #4096 r268 = ~r268;
  always #8192 r269 = ~r269;
  always #16384 r270 = ~r270;
  always #32768 r271 = ~r271;
  always #65536 r272 = ~r272;
  always #131072 r273 = ~r273;
  always #262144 r274 = ~r274;
  always #524288 r275 = ~r275;
  always #1048576 r276 = ~r276;
  always #2097152 r277 = ~r277;
  always #4194304 r278 = ~r278;
  always #8388608 r279 = ~r279;
  always #16777216 r280 = ~r280;
  always #33554432 r281 = ~r281;
  always #67108864 r282 = ~r282;
  always #134217728 r283 = ~r283;
  always #268435456 r284 = ~r284;
  always #536870912 r285 = ~r285;
  always #1073741824 r286 = ~r286;
  always #2147483648 r287 = ~r287;
  always #4294967296 r288 = ~r288;
  always #8589934592 r289 = ~r289;
  always #17179869184 r290 = ~r290;
  always #34359738368 r291 = ~r291;
  always #68719476736 r292 = ~r292;
  always #137438953472 r293 = ~r293;
  always #274877906944 r294 = ~r294;
  always #549755813888 r295 = ~r295;
  always #1099511627776 r296 = ~r296;
  always #2199023255552 r297 = ~r297;
  always #4398046511104 r298 = ~r298;
  always #8796093022208 r299 = ~r299;
  always #17592186044416 r300 = ~r300;
  always #35184372088832 r301 = ~r301;
  always #70368744177664 r302 = ~r302;
  always #140737488355328 r303 = ~r303;
  always #281474976710656 r304 = ~r304;
  always #562949953421312 r305 = ~r305;
  always #1125899906842624 r306 = ~r306;
  always #2251799813685248 r307 = ~r307;
  always #4503599627370496 r308 = ~r308;
  always #9007199254740992 r309 = ~r309;
  always #18014398509481984 r310 = ~r310;
  always #36028797018963968 r311 = ~r311;
  always #72057594037927936 r312 = ~r312;
  always #144115188075855872 r313 = ~r313;
  always #288230376151711744 r314 = ~r314;
  always #576460752303423488 r315 = ~r315;
  always #1152921504606846976 r316 = ~r316;
  always #2305843009213693952 r317 = ~r317;
  always #4611686018427387904 r318 = ~r318;
  always #9223372036854775808 r319 = ~r319;
  always #1 r320 = ~r320;
  always #2 r321 = ~r321;
  always #4 r322 = ~r322;
  always #8 r323 = ~r323;
  always #16 r324 = ~r324;
  always #32 r325 = ~r325;
  always #64 r326 = ~r326;
  always #128 r327 = ~r327;
  always #256 r328 = ~r328;
  always #512 r329 = ~r329;
  always #1024 r330 = ~r330;
  always #2048 r331 = ~r331;
  always #4096 r332 = ~r332;
  always #8192 r333 = ~r333;
  always #16384 r334 = ~r334;
  always #32768 r335 = ~r335;
  always #65536 r336 = ~r336;
  always #131072 r337 = ~r337;
  always #262144 r338 = ~r338;
  always #524288 r339 = ~r339;
  always #1048576 r340 = ~r340;
  always #2097152 r341 = ~r341;
  always #4194304 r342 = ~r342;
  always #8388608 r343 = ~r343;
  always #16777216 r344 = ~r344;
  always #33554432 r345 = ~r345;
  always #67108864 r346 = ~r346;
  always #134217728 r347 = ~r347;
  always #268435456 r348 = ~r348;
  always #536870912 r349 = ~r349;
  always #1073741824 r350 = ~r350;
  always #2147483648 r351 = ~r351;
  always #4294967296 r352 = ~r352;
  always #8589934592 r353 = ~r353;
  always #17179869184 r354 = ~r354;
  always #34359738368 r355 = ~r355;
  always #68719476736 r356 = ~r356;
  always #137438953472 r357 = ~r357;
  always #274877906944 r358 = ~r358;
  always #549755813888 r359 = ~r359;
  always #1099511627776 r360 = ~r360;
  always #2199023255552 r361 = ~r361;
  always #4398046511104 r362 = ~r362;
  always #8796093022208 r363 = ~r363;
  always #17592186044416 r364 = ~r364;
  always #35184372088832 r365 = ~r365;
  always #70368744177664 r366 = ~r366;
  always #140737488355328 r367 = ~r367;
  always #281474976710656 r368 = ~r368;
  always #562949953421312 r369 = ~r369;
  always #1125899906842624 r370 = ~r370;
  always #2251799813685248 r371 = ~r371;
  always #4503599627370496 r372 = ~r372;
  always #9007199254740992 r373 = ~r373;
  always #18014398509481984 r374 = ~r374;
  always #36028797018963968 r375 = ~r375;
  always #72057594037927936 r376 = ~r376;
  always #144115188075855872 r377 = ~r377;
  always #288230376151711744 r378 = ~r378;
  always #576460752303423488 r379 = ~r379;
  always #1152921504606846976 r380 = ~r380;
  always #2305843009213693952 r381 = ~r381;
  always #4611686018427387904 r382 = ~r382;
  always #9223372036854775808 r383 = ~r383;
  always #1 r384 = ~r384;
  always #2 r385 = ~r385;
  always #4 r386 = ~r386;
  always #8 r387 = ~r387;
  always #16 r388 = ~r388;
  always #32 r389 = ~r389;
  always #64 r390 = ~r390;
  always #128 r391 = ~r391;
  always #256 r392 = ~r392;
  always #512 r393 = ~r393;
  always #1024 r394 = ~r394;
  always #2048 r395 = ~r395;
  always #4096 r396 = ~r396;
  always #8192 r397 = ~r397;
  always #16384 r398 = ~r398;
  always #32768 r399 = ~r399;
  always #65536 r400 = ~r400;
  always #131072 r401 = ~r401;
  always #262144 r402 = ~r402;
  always #524288 r403 = ~r403;
  always #1048576 r404 = ~r404;
  always #2097152 r405 = ~r405;
  always #4194304 r406 = ~r406;
  always #8388608 r407 = ~r407;
  always #16777216 r408 = ~r408;
  always #33554432 r409 = ~r409;
  always #67108864 r410 = ~r410;
  always #134217728 r411 = ~r411;
  always #268435456 r412 = ~r412;
  always #536870912 r413 = ~r413;
  always #1073741824 r414 = ~r414;
  always #2147483648 r415 = ~r415;
  always #4294967296 r416 = ~r416;
  always #8589934592 r417 = ~r417;
  always #17179869184 r418 = ~r418;
  always #34359738368 r419 = ~r419;
  always #68719476736 r420 = ~r420;
  always #137438953472 r421 = ~r421;
  always #274877906944 r422 = ~r422;
  always #549755813888 r423 = ~r423;
  always #1099511627776 r424 = ~r424;
  always #2199023255552 r425 = ~r425;
  always #4398046511104 r426 = ~r426;
  always #8796093022208 r427 = ~r427;
  always #17592186044416 r428 = ~r428;
  always #35184372088832 r429 = ~r429;
  always #70368744177664 r430 = ~r430;
  always #140737488355328 r431 = ~r431;
  always #281474976710656 r432 = ~r432;
  always #562949953421312 r433 = ~r433;
  always #1125899906842624 r434 = ~r434;
  always #2251799813685248 r435 = ~r435;
  always #4503599627370496 r436 = ~r436;
  always #9007199254740992 r437 = ~r437;
  always #18014398509481984 r438 = ~r438;
  always #36028797018963968 r439 = ~r439;
  always #72057594037927936 r440 = ~r440;
  always #144115188075855872 r441 = ~r441;
  always #288230376151711744 r442 = ~r442;
  always #576460752303423488 r443 = ~r443;
  always #1152921504606846976 r444 = ~r444;
  always #2305843009213693952 r445 = ~r445;
  always #4611686018427387904 r446 = ~r446;
  always #9223372036854775808 r447 = ~r447;
  always #1 r448 = ~r448;
  always #2 r449 = ~r449;
  always #4 r450 = ~r450;
  always #8 r451 = ~r451;
  always #16 r452 = ~r452;
  always #32 r453 = ~r453;
  always #64 r454 = ~r454;
  always #128 r455 = ~r455;
  always #256 r456 = ~r456;
  always #512 r457 = ~r457;
  always #1024 r458 = ~r458;
  always #2048 r459 = ~r459;
  always #4096 r460 = ~r460;
  always #8192 r461 = ~r461;
  always #16384 r462 = ~r462;
  always #32768 r463 = ~r463;
  always #65536 r464 = ~r464;
  always #131072 r465 = ~r465;
  always #262144 r466 = ~r466;
  always #524288 r467 = ~r467;
  always #1048576 r468 = ~r468;
  always #2097152 r469 = ~r469;
  always #4194304 r470 = ~r470;
  always #8388608 r471 = ~r471;
  always #16777216 r472 = ~r472;
  always #33554432 r473 = ~r473;
  always #67108864 r474 = ~r474;
  always #134217728 r475 = ~r475;
  always #268435456 r476 = ~r476;
  always #536870912 r477 = ~r477;
  always #1073741824 r478 = ~r478;
  always #2147483648 r479 = ~r479;
  always #4294967296 r480 = ~r480;
  always #8589934592 r481 = ~r481;
  always #17179869184 r482 = ~r482;
  always #34359738368 r483 = ~r483;
  always #68719476736 r484 = ~r484;
  always #137438953472 r485 = ~r485;
  always #274877906944 r486 = ~r486;
  always #549755813888 r487 = ~r487;
  always #1099511627776 r488 = ~r488;
  always #2199023255552 r489 = ~r489;
  always #4398046511104 r490 = ~r490;
  always #8796093022208 r491 = ~r491;
  always #17592186044416 r492 = ~r492;
  always #35184372088832 r493 = ~r493;
  always #70368744177664 r494 = ~r494;
  always #140737488355328 r495 = ~r495;
  always #281474976710656 r496 = ~r496;
endmodule
*/
// ****** TestBench Module Defination End ******

/*
// ******* The results for this case *********
******* result_1.txt *********
1)
  Loop Signals: w_139_229, w_139_230, w_139_231, 
  Loop Gates: I139_228.port2, I139_229.port2, I139_230.port2, 

2)
  Loop Signals: w_489_323, w_489_324, w_489_325, w_489_326, w_489_327, w_489_328, w_489_329, w_489_330, w_489_331, w_489_332, 
  Loop Gates: I489_322.port1, I489_323.port2, I489_324.port1, I489_325.port1, I489_326.port2, I489_327.port1, I489_328.port1, I489_329.port1, I489_330.port1, I489_331.port1, 

3)
  Loop Signals: w_489_325, w_489_336, w_489_337, w_489_338, w_489_339, w_489_340, w_489_341, w_489_342, w_489_344, 
  Loop Gates: I489_323.port1, I489_332.port1, I489_333.port1, I489_334.port1, I489_335.port2, I489_336.port1, I489_337.port1, I489_338.port1, I489_339.port2, 

4)
  Loop Signals: w_158_038, w_158_039, w_158_040, w_158_041, w_158_042, w_158_043, w_158_044, w_158_045, w_158_046, w_158_047, w_158_048, 
  Loop Gates: I158_037.port2, I158_038.port1, I158_039.port1, I158_040.port1, I158_041.port1, I158_042.port1, I158_043.port2, I158_044.port1, I158_045.port1, I158_046.port1, I158_047.port2, 

5)
  Loop Signals: w_431_274, w_431_275, w_431_276, w_431_277, 
  Loop Gates: I431_273.port2, I431_274.port1, I431_275.port2, I431_276.port2, 

6)
  Loop Signals: w_431_275, w_431_281, w_431_282, w_431_283, w_431_284, w_431_285, w_431_286, w_431_287, w_431_288, w_431_290, 
  Loop Gates: I431_273.port1, I431_277.port2, I431_278.port1, I431_279.port1, I431_280.port1, I431_281.port1, I431_282.port2, I431_283.port1, I431_284.port1, I431_285.port2, 

7)
  Loop Signals: w_029_249, w_029_250, w_029_251, w_029_252, w_029_253, w_029_254, w_029_255, w_029_256, 
  Loop Gates: I029_248.port2, I029_249.port1, I029_250.port1, I029_251.port1, I029_252.port1, I029_253.port1, I029_254.port1, I029_255.port2, 

8)
  Loop Signals: w_029_256, w_029_260, w_029_261, w_029_262, w_029_263, w_029_265, 
  Loop Gates: I029_254.port2, I029_256.port2, I029_257.port2, I029_258.port2, I029_259.port1, I029_260.port2, 

9)
  Loop Signals: w_082_340, w_082_341, w_082_342, w_082_343, w_082_344, w_082_345, 
  Loop Gates: I082_339.port2, I082_340.port1, I082_341.port1, I082_342.port1, I082_343.port1, I082_344.port2, 

10)
  Loop Signals: w_445_400, w_445_401, w_445_402, w_445_403, w_445_404, 
  Loop Gates: I445_399.port1, I445_400.port1, I445_401.port2, I445_402.port2, I445_403.port1, 

11)
  Loop Signals: w_445_402, w_445_408, w_445_409, w_445_410, w_445_411, w_445_412, w_445_413, w_445_414, w_445_416, 
  Loop Gates: I445_400.port2, I445_404.port2, I445_405.port1, I445_406.port1, I445_407.port2, I445_408.port2, I445_409.port2, I445_410.port1, I445_411.port2, 

12)
  Loop Signals: w_285_025, w_285_026, w_285_027, w_285_028, w_285_029, w_285_030, w_285_031, w_285_032, w_285_033, w_285_034, w_285_035, 
  Loop Gates: I285_024.port1, I285_025.port1, I285_026.port1, I285_027.port1, I285_028.port2, I285_029.port1, I285_030.port1, I285_031.port2, I285_032.port2, I285_033.port1, I285_034.port2, 

13)
  Loop Signals: w_186_061, w_186_062, w_186_063, w_186_064, w_186_065, w_186_066, w_186_067, w_186_068, 
  Loop Gates: I186_060.port1, I186_061.port1, I186_062.port1, I186_063.port1, I186_064.port2, I186_065.port2, I186_066.port1, I186_067.port1, 

14)
  Loop Signals: w_186_065, w_186_072, w_186_073, w_186_074, w_186_075, w_186_076, w_186_077, w_186_078, w_186_079, w_186_080, w_186_081, w_186_082, w_186_083, w_186_085, 
  Loop Gates: I186_063.port2, I186_068.port1, I186_069.port2, I186_070.port2, I186_071.port2, I186_072.port1, I186_073.port1, I186_074.port2, I186_075.port1, I186_076.port2, I186_077.port1, I186_078.port2, I186_079.port1, I186_080.port2, 

15)
  Loop Signals: w_338_357, w_338_358, w_338_359, w_338_360, w_338_361, w_338_362, 
  Loop Gates: I338_356.port2, I338_357.port1, I338_358.port2, I338_359.port2, I338_360.port1, I338_361.port1, 

16)
  Loop Signals: w_088_454, w_088_455, w_088_456, 
  Loop Gates: I088_453.port1, I088_454.port1, I088_455.port1, 

17)
  Loop Signals: w_088_456, w_088_460, w_088_461, w_088_462, w_088_463, w_088_464, w_088_465, w_088_466, w_088_467, w_088_468, w_088_469, w_088_471, 
  Loop Gates: I088_454.port2, I088_456.port2, I088_457.port2, I088_458.port2, I088_459.port1, I088_460.port2, I088_461.port1, I088_462.port1, I088_463.port1, I088_464.port2, I088_465.port1, I088_466.port2, 

18)
  Loop Signals: w_372_147, w_372_148, w_372_149, w_372_150, w_372_151, w_372_152, w_372_153, w_372_154, 
  Loop Gates: I372_146.port1, I372_147.port1, I372_148.port1, I372_149.port2, I372_150.port2, I372_151.port1, I372_152.port1, I372_153.port1, 

19)
  Loop Signals: w_484_092, w_484_093, w_484_094, w_484_095, w_484_096, 
  Loop Gates: I484_091.port1, I484_092.port1, I484_093.port1, I484_094.port1, I484_095.port1, 

20)
  Loop Signals: w_484_096, w_484_100, w_484_101, w_484_102, w_484_103, w_484_105, 
  Loop Gates: I484_094.port2, I484_096.port1, I484_097.port1, I484_098.port1, I484_099.port1, I484_100.port2, 

21)
  Loop Signals: w_203_367, w_203_368, w_203_369, w_203_370, w_203_371, w_203_372, w_203_373, 
  Loop Gates: I203_366.port1, I203_367.port2, I203_368.port1, I203_369.port1, I203_370.port2, I203_371.port1, I203_372.port1, 

22)
  Loop Signals: w_203_369, w_203_377, w_203_378, w_203_379, w_203_380, w_203_381, w_203_382, w_203_383, w_203_384, w_203_385, w_203_386, w_203_387, w_203_388, w_203_390, 
  Loop Gates: I203_367.port1, I203_373.port1, I203_374.port1, I203_375.port1, I203_376.port1, I203_377.port1, I203_378.port1, I203_379.port1, I203_380.port1, I203_381.port1, I203_382.port1, I203_383.port2, I203_384.port1, I203_385.port2, 

23)
  Loop Signals: w_476_252, w_476_253, w_476_254, w_476_255, w_476_256, w_476_257, w_476_258, w_476_259, w_476_260, 
  Loop Gates: I476_251.port1, I476_252.port1, I476_253.port1, I476_254.port2, I476_255.port1, I476_256.port1, I476_257.port1, I476_258.port2, I476_259.port2, 

24)
  Loop Signals: w_138_241, w_138_242, w_138_243, w_138_244, w_138_245, w_138_246, w_138_247, w_138_248, 
  Loop Gates: I138_240.port1, I138_241.port2, I138_242.port2, I138_243.port1, I138_244.port1, I138_245.port1, I138_246.port1, I138_247.port1, 

25)
  Loop Signals: w_138_244, w_138_252, w_138_253, w_138_254, w_138_255, w_138_256, w_138_257, w_138_259, 
  Loop Gates: I138_242.port1, I138_248.port1, I138_249.port2, I138_250.port2, I138_251.port1, I138_252.port1, I138_253.port1, I138_254.port2, 

26)
  Loop Signals: w_373_102, w_373_103, w_373_104, w_373_105, w_373_106, w_373_107, 
  Loop Gates: I373_102.port1, I373_103.port2, I373_104.port1, I373_105.port2, I373_106.port2, I373_107.port1, 

27)
  Loop Signals: w_127_492, w_127_493, w_127_494, w_127_495, w_127_496, w_127_497, w_127_498, w_127_499, w_127_500, w_127_501, w_127_502, w_127_503, 
  Loop Gates: I127_491.port1, I127_492.port1, I127_493.port1, I127_494.port1, I127_495.port1, I127_496.port1, I127_497.port1, I127_498.port1, I127_499.port1, I127_500.port1, I127_501.port1, I127_502.port1, 

28)
  Loop Signals: w_487_077, w_487_078, w_487_079, 
  Loop Gates: I487_076.port1, I487_077.port2, I487_078.port1, 

29)
  Loop Signals: w_487_077, w_487_083, w_487_084, w_487_085, w_487_086, w_487_087, w_487_088, w_487_089, w_487_090, w_487_091, w_487_092, w_487_093, w_487_094, w_487_096, 
  Loop Gates: I487_078.port2, I487_079.port1, I487_080.port1, I487_081.port2, I487_082.port2, I487_083.port1, I487_084.port2, I487_085.port2, I487_086.port2, I487_087.port2, I487_088.port2, I487_089.port1, I487_090.port1, I487_091.port2, 

30)
  Loop Signals: w_039_499, w_039_500, w_039_501, w_039_502, w_039_503, w_039_504, w_039_505, w_039_506, w_039_507, w_039_508, w_039_509, 
  Loop Gates: I039_498.port1, I039_499.port1, I039_500.port1, I039_501.port2, I039_502.port2, I039_503.port1, I039_504.port1, I039_505.port2, I039_506.port1, I039_507.port1, I039_508.port2, 

31)
  Loop Signals: w_039_500, w_039_513, w_039_514, w_039_515, w_039_516, w_039_517, w_039_518, w_039_519, w_039_520, w_039_522, 
  Loop Gates: I039_498.port2, I039_509.port1, I039_510.port2, I039_511.port1, I039_512.port1, I039_513.port1, I039_514.port2, I039_515.port1, I039_516.port1, I039_517.port2, 

32)
  Loop Signals: w_114_266, w_114_267, w_114_268, w_114_269, w_114_270, w_114_271, w_114_272, w_114_273, w_114_274, w_114_275, w_114_276, 
  Loop Gates: I114_265.port1, I114_266.port1, I114_267.port1, I114_268.port1, I114_269.port2, I114_270.port2, I114_271.port1, I114_272.port2, I114_273.port2, I114_274.port2, I114_275.port2, 

33)
  Loop Signals: w_114_276, w_114_280, w_114_281, w_114_282, w_114_283, w_114_284, w_114_285, w_114_286, w_114_287, w_114_289, 
  Loop Gates: I114_274.port1, I114_276.port1, I114_277.port2, I114_278.port2, I114_279.port1, I114_280.port2, I114_281.port1, I114_282.port2, I114_283.port1, I114_284.port2, 

34)
  Loop Signals: w_192_260, w_192_261, w_192_262, w_192_263, w_192_264, w_192_265, w_192_266, w_192_267, w_192_268, 
  Loop Gates: I192_259.port1, I192_260.port1, I192_261.port2, I192_262.port1, I192_263.port2, I192_264.port1, I192_265.port1, I192_266.port2, I192_267.port1, 

35)
  Loop Signals: w_226_396, w_226_397, w_226_398, w_226_399, w_226_400, w_226_401, w_226_402, w_226_403, 
  Loop Gates: I226_395.port1, I226_396.port1, I226_397.port2, I226_398.port1, I226_399.port1, I226_400.port1, I226_401.port1, I226_402.port1, 

36)
  Loop Signals: w_317_341, w_317_342, w_317_343, w_317_344, w_317_345, w_317_346, w_317_347, w_317_348, w_317_349, w_317_350, w_317_351, 
  Loop Gates: I317_340.port2, I317_341.port1, I317_342.port1, I317_343.port1, I317_344.port2, I317_345.port2, I317_346.port1, I317_347.port1, I317_348.port2, I317_349.port1, I317_350.port1, 

37)
  Loop Signals: w_303_197, w_303_198, w_303_199, w_303_200, 
  Loop Gates: I303_196.port2, I303_197.port1, I303_198.port2, I303_199.port1, 

38)
  Loop Signals: w_303_198, w_303_204, w_303_205, w_303_206, w_303_207, w_303_208, w_303_209, w_303_210, w_303_211, w_303_212, w_303_213, w_303_215, 
  Loop Gates: I303_196.port1, I303_200.port1, I303_201.port1, I303_202.port1, I303_203.port1, I303_204.port1, I303_205.port1, I303_206.port1, I303_207.port2, I303_208.port1, I303_209.port1, I303_210.port2, 

39)
  Loop Signals: w_318_382, w_318_383, w_318_384, w_318_385, w_318_386, w_318_387, w_318_388, w_318_389, w_318_390, 
  Loop Gates: I318_382.port1, I318_383.port1, I318_384.port1, I318_385.port2, I318_386.port1, I318_387.port1, I318_388.port1, I318_389.port2, I318_390.port1, 

40)
  Loop Signals: w_318_385, w_318_394, w_318_395, w_318_396, w_318_397, w_318_398, w_318_399, w_318_401, 
  Loop Gates: I318_384.port2, I318_391.port2, I318_392.port1, I318_393.port1, I318_394.port2, I318_395.port1, I318_396.port1, I318_397.port2, 

41)
  Loop Signals: w_375_263, w_375_264, w_375_265, w_375_266, w_375_267, w_375_268, w_375_269, w_375_270, w_375_271, w_375_272, 
  Loop Gates: I375_262.port1, I375_263.port1, I375_264.port1, I375_265.port2, I375_266.port2, I375_267.port1, I375_268.port1, I375_269.port1, I375_270.port1, I375_271.port1, 

42)
  Loop Signals: w_375_267, w_375_276, w_375_277, w_375_278, w_375_279, w_375_280, w_375_281, w_375_282, w_375_283, w_375_284, w_375_285, w_375_286, w_375_288, 
  Loop Gates: I375_265.port1, I375_272.port2, I375_273.port1, I375_274.port2, I375_275.port1, I375_276.port2, I375_277.port2, I375_278.port1, I375_279.port1, I375_280.port2, I375_281.port2, I375_282.port1, I375_283.port2, 

43)
  Loop Signals: w_262_063, w_262_064, w_262_065, w_262_066, w_262_067, w_262_068, w_262_069, w_262_070, w_262_071, w_262_072, w_262_073, w_262_074, 
  Loop Gates: I262_062.port1, I262_063.port2, I262_064.port2, I262_065.port2, I262_066.port1, I262_067.port1, I262_068.port1, I262_069.port2, I262_070.port1, I262_071.port1, I262_072.port2, I262_073.port2, 

44)
  Loop Signals: w_093_426, w_093_427, w_093_428, w_093_429, w_093_430, 
  Loop Gates: I093_425.port1, I093_426.port1, I093_427.port2, I093_428.port1, I093_429.port2, 

45)
  Loop Signals: w_093_429, w_093_434, w_093_435, w_093_436, w_093_437, w_093_438, w_093_439, w_093_440, w_093_441, w_093_442, w_093_443, w_093_444, w_093_445, w_093_447, 
  Loop Gates: I093_427.port1, I093_430.port1, I093_431.port1, I093_432.port1, I093_433.port1, I093_434.port2, I093_435.port2, I093_436.port1, I093_437.port1, I093_438.port2, I093_439.port2, I093_440.port1, I093_441.port1, I093_442.port2, 

46)
  Loop Signals: w_127_507, w_127_508, w_127_509, w_127_510, w_127_511, w_127_512, w_127_513, w_127_514, w_127_515, w_127_516, w_127_517, 
  Loop Gates: I127_503.port2, I127_504.port2, I127_505.port1, I127_506.port2, I127_507.port2, I127_508.port2, I127_509.port1, I127_510.port2, I127_511.port2, I127_512.port1, I127_513.port1, 

47)
  Loop Signals: w_127_515, w_127_521, w_127_522, w_127_523, w_127_524, w_127_525, w_127_526, w_127_527, w_127_528, w_127_529, w_127_530, w_127_531, w_127_532, w_127_534, 
  Loop Gates: I127_510.port1, I127_514.port1, I127_515.port1, I127_516.port1, I127_517.port1, I127_518.port2, I127_519.port2, I127_520.port2, I127_521.port1, I127_522.port1, I127_523.port2, I127_524.port1, I127_525.port1, I127_526.port2, 

48)
  Loop Signals: w_022_164, w_022_165, w_022_166, w_022_167, w_022_168, w_022_169, w_022_170, w_022_171, w_022_172, w_022_173, 
  Loop Gates: I022_163.port2, I022_164.port1, I022_165.port1, I022_166.port1, I022_167.port2, I022_168.port2, I022_169.port1, I022_170.port2, I022_171.port2, I022_172.port2, 

49)
  Loop Signals: w_164_188, w_164_189, w_164_190, w_164_191, w_164_192, w_164_193, w_164_194, w_164_195, 
  Loop Gates: I164_187.port1, I164_188.port1, I164_189.port2, I164_190.port1, I164_191.port2, I164_192.port2, I164_193.port1, I164_194.port1, 

50)
  Loop Signals: w_173_283, w_173_284, w_173_285, w_173_286, w_173_287, w_173_288, w_173_289, w_173_290, w_173_291, w_173_292, 
  Loop Gates: I173_282.port1, I173_283.port1, I173_284.port2, I173_285.port2, I173_286.port1, I173_287.port2, I173_288.port1, I173_289.port2, I173_290.port1, I173_291.port2, 

******* result_2.txt *********
1)
  Loop Signals: w_489_323, w_489_324, w_489_325, w_489_326, w_489_327, w_489_328, w_489_329, w_489_330, w_489_331, w_489_332, 
  Loop Gates: I489_322.port1, I489_323.port2, I489_324.port1, I489_325.port1, I489_326.port2, I489_327.port1, I489_328.port1, I489_329.port1, I489_330.port1, I489_331.port1, 

2)
  Loop Signals: w_431_275, w_431_281, w_431_282, w_431_283, w_431_284, w_431_285, w_431_286, w_431_287, w_431_288, w_431_290, 
  Loop Gates: I431_273.port1, I431_277.port2, I431_278.port1, I431_279.port1, I431_280.port1, I431_281.port1, I431_282.port2, I431_283.port1, I431_284.port1, I431_285.port2, 

3)
  Loop Signals: w_029_249, w_029_250, w_029_251, w_029_252, w_029_253, w_029_254, w_029_255, w_029_256, 
  Loop Gates: I029_248.port2, I029_249.port1, I029_250.port1, I029_251.port1, I029_252.port1, I029_253.port1, I029_254.port1, I029_255.port2, 

4)
  Loop Signals: w_285_025, w_285_026, w_285_027, w_285_028, w_285_029, w_285_030, w_285_031, w_285_032, w_285_033, w_285_034, w_285_035, 
  Loop Gates: I285_024.port1, I285_025.port1, I285_026.port1, I285_027.port1, I285_028.port2, I285_029.port1, I285_030.port1, I285_031.port2, I285_032.port2, I285_033.port1, I285_034.port2, 

5)
  Loop Signals: w_338_357, w_338_358, w_338_359, w_338_360, w_338_361, w_338_362, 
  Loop Gates: I338_356.port2, I338_357.port1, I338_358.port2, I338_359.port2, I338_360.port1, I338_361.port1, 

6)
  Loop Signals: w_088_454, w_088_455, w_088_456, 
  Loop Gates: I088_453.port1, I088_454.port1, I088_455.port1, 

7)
  Loop Signals: w_484_096, w_484_100, w_484_101, w_484_102, w_484_103, w_484_105, 
  Loop Gates: I484_094.port2, I484_096.port1, I484_097.port1, I484_098.port1, I484_099.port1, I484_100.port2, 

8)
  Loop Signals: w_203_369, w_203_377, w_203_378, w_203_379, w_203_380, w_203_381, w_203_382, w_203_383, w_203_384, w_203_385, w_203_386, w_203_387, w_203_388, w_203_390, 
  Loop Gates: I203_367.port1, I203_373.port1, I203_374.port1, I203_375.port1, I203_376.port1, I203_377.port1, I203_378.port1, I203_379.port1, I203_380.port1, I203_381.port1, I203_382.port1, I203_383.port2, I203_384.port1, I203_385.port2, 

9)
  Loop Signals: w_476_252, w_476_253, w_476_254, w_476_255, w_476_256, w_476_257, w_476_258, w_476_259, w_476_260, 
  Loop Gates: I476_251.port1, I476_252.port1, I476_253.port1, I476_254.port2, I476_255.port1, I476_256.port1, I476_257.port1, I476_258.port2, I476_259.port2, 

10)
  Loop Signals: w_373_102, w_373_103, w_373_104, w_373_105, w_373_106, w_373_107, 
  Loop Gates: I373_102.port1, I373_103.port2, I373_104.port1, I373_105.port2, I373_106.port2, I373_107.port1, 

11)
  Loop Signals: w_127_492, w_127_493, w_127_494, w_127_495, w_127_496, w_127_497, w_127_498, w_127_499, w_127_500, w_127_501, w_127_502, w_127_503, 
  Loop Gates: I127_491.port1, I127_492.port1, I127_493.port1, I127_494.port1, I127_495.port1, I127_496.port1, I127_497.port1, I127_498.port1, I127_499.port1, I127_500.port1, I127_501.port1, I127_502.port1, 

12)
  Loop Signals: w_487_077, w_487_078, w_487_079, 
  Loop Gates: I487_076.port1, I487_077.port2, I487_078.port1, 

13)
  Loop Signals: w_487_077, w_487_083, w_487_084, w_487_085, w_487_086, w_487_087, w_487_088, w_487_089, w_487_090, w_487_091, w_487_092, w_487_093, w_487_094, w_487_096, 
  Loop Gates: I487_078.port2, I487_079.port1, I487_080.port1, I487_081.port2, I487_082.port2, I487_083.port1, I487_084.port2, I487_085.port2, I487_086.port2, I487_087.port2, I487_088.port2, I487_089.port1, I487_090.port1, I487_091.port2, 

14)
  Loop Signals: w_039_499, w_039_500, w_039_501, w_039_502, w_039_503, w_039_504, w_039_505, w_039_506, w_039_507, w_039_508, w_039_509, 
  Loop Gates: I039_498.port1, I039_499.port1, I039_500.port1, I039_501.port2, I039_502.port2, I039_503.port1, I039_504.port1, I039_505.port2, I039_506.port1, I039_507.port1, I039_508.port2, 

15)
  Loop Signals: w_114_266, w_114_267, w_114_268, w_114_269, w_114_270, w_114_271, w_114_272, w_114_273, w_114_274, w_114_275, w_114_276, 
  Loop Gates: I114_265.port1, I114_266.port1, I114_267.port1, I114_268.port1, I114_269.port2, I114_270.port2, I114_271.port1, I114_272.port2, I114_273.port2, I114_274.port2, I114_275.port2, 

16)
  Loop Signals: w_114_276, w_114_280, w_114_281, w_114_282, w_114_283, w_114_284, w_114_285, w_114_286, w_114_287, w_114_289, 
  Loop Gates: I114_274.port1, I114_276.port1, I114_277.port2, I114_278.port2, I114_279.port1, I114_280.port2, I114_281.port1, I114_282.port2, I114_283.port1, I114_284.port2, 

17)
  Loop Signals: w_192_260, w_192_261, w_192_262, w_192_263, w_192_264, w_192_265, w_192_266, w_192_267, w_192_268, 
  Loop Gates: I192_259.port1, I192_260.port1, I192_261.port2, I192_262.port1, I192_263.port2, I192_264.port1, I192_265.port1, I192_266.port2, I192_267.port1, 

18)
  Loop Signals: w_318_382, w_318_383, w_318_384, w_318_385, w_318_386, w_318_387, w_318_388, w_318_389, w_318_390, 
  Loop Gates: I318_382.port1, I318_383.port1, I318_384.port1, I318_385.port2, I318_386.port1, I318_387.port1, I318_388.port1, I318_389.port2, I318_390.port1, 

19)
  Loop Signals: w_375_263, w_375_264, w_375_265, w_375_266, w_375_267, w_375_268, w_375_269, w_375_270, w_375_271, w_375_272, 
  Loop Gates: I375_262.port1, I375_263.port1, I375_264.port1, I375_265.port2, I375_266.port2, I375_267.port1, I375_268.port1, I375_269.port1, I375_270.port1, I375_271.port1, 

20)
  Loop Signals: w_262_063, w_262_064, w_262_065, w_262_066, w_262_067, w_262_068, w_262_069, w_262_070, w_262_071, w_262_072, w_262_073, w_262_074, 
  Loop Gates: I262_062.port1, I262_063.port2, I262_064.port2, I262_065.port2, I262_066.port1, I262_067.port1, I262_068.port1, I262_069.port2, I262_070.port1, I262_071.port1, I262_072.port2, I262_073.port2, 

21)
  Loop Signals: w_093_426, w_093_427, w_093_428, w_093_429, w_093_430, 
  Loop Gates: I093_425.port1, I093_426.port1, I093_427.port2, I093_428.port1, I093_429.port2, 

22)
  Loop Signals: w_127_515, w_127_521, w_127_522, w_127_523, w_127_524, w_127_525, w_127_526, w_127_527, w_127_528, w_127_529, w_127_530, w_127_531, w_127_532, w_127_534, 
  Loop Gates: I127_510.port1, I127_514.port1, I127_515.port1, I127_516.port1, I127_517.port1, I127_518.port2, I127_519.port2, I127_520.port2, I127_521.port1, I127_522.port1, I127_523.port2, I127_524.port1, I127_525.port1, I127_526.port2, 

23)
  Loop Signals: w_164_188, w_164_189, w_164_190, w_164_191, w_164_192, w_164_193, w_164_194, w_164_195, 
  Loop Gates: I164_187.port1, I164_188.port1, I164_189.port2, I164_190.port1, I164_191.port2, I164_192.port2, I164_193.port1, I164_194.port1, 

******* result_3.txt *********
1)
  Loop Signals: w_139_229, w_139_230, w_139_231, 
  Loop Gates: I139_228.port2, I139_229.port2, I139_230.port2, 
  Loop Conditions: I139_228.port1=1, I139_229.port1=0, I139_230.port1=1, 
  (Singal Values: w_044_133=1, w_070_095=1, w_112_232=0, )

2)
  Loop Signals: w_489_325, w_489_336, w_489_337, w_489_338, w_489_339, w_489_340, w_489_341, w_489_342, w_489_344, 
  Loop Gates: I489_323.port1, I489_332.port1, I489_333.port1, I489_334.port1, I489_335.port2, I489_336.port1, I489_337.port1, I489_338.port1, I489_339.port2, 
  Loop Conditions: I489_323.port2=0, I489_332.port2=0, I489_333.port2=1, I489_334.port2=1, I489_335.port1=0, I489_337.port2=1, I489_339.port1=1, 
  (Singal Values: w_069_069=0, w_187_131=1, w_244_089=0, w_405_178=1, w_413_052=1, w_423_096=1, w_489_324=0, )

3)
  Loop Signals: w_158_038, w_158_039, w_158_040, w_158_041, w_158_042, w_158_043, w_158_044, w_158_045, w_158_046, w_158_047, w_158_048, 
  Loop Gates: I158_037.port2, I158_038.port1, I158_039.port1, I158_040.port1, I158_041.port1, I158_042.port1, I158_043.port2, I158_044.port1, I158_045.port1, I158_046.port1, I158_047.port2, 
  Loop Conditions: I158_037.port1=0, I158_038.port2=1, I158_040.port2=1, I158_041.port2=1, I158_042.port2=1, I158_043.port1=0, I158_044.port2=1, I158_045.port2=1, I158_047.port1=0, 
  (Singal Values: w_005_219=0, w_006_000=1, w_057_036=0, w_074_004=1, w_075_124=1, w_101_039=1, w_127_260=1, w_129_000=0, w_147_127=1, )

4)
  Loop Signals: w_431_274, w_431_275, w_431_276, w_431_277, 
  Loop Gates: I431_273.port2, I431_274.port1, I431_275.port2, I431_276.port2, 
  Loop Conditions: I431_273.port1=0, I431_275.port1=0, I431_276.port1=0, 
  (Singal Values: w_016_118=0, w_249_102=0, w_431_290=0, )

5)
  Loop Signals: w_029_256, w_029_260, w_029_261, w_029_262, w_029_263, w_029_265, 
  Loop Gates: I029_254.port2, I029_256.port2, I029_257.port2, I029_258.port2, I029_259.port1, I029_260.port2, 
  Loop Conditions: I029_254.port1=1, I029_256.port1=0, I029_257.port1=0, I029_258.port1=0, I029_260.port1=1, 
  (Singal Values: w_003_069=0, w_020_055=1, w_022_131=0, w_028_085=0, w_029_255=1, )

6)
  Loop Signals: w_082_340, w_082_341, w_082_342, w_082_343, w_082_344, w_082_345, 
  Loop Gates: I082_339.port2, I082_340.port1, I082_341.port1, I082_342.port1, I082_343.port1, I082_344.port2, 
  Loop Conditions: I082_339.port1=1, I082_340.port2=0, I082_342.port2=0, I082_344.port1=1, 
  (Singal Values: w_007_357=1, w_017_104=0, w_057_048=0, w_080_021=1, )

7)
  Loop Signals: w_445_400, w_445_401, w_445_402, w_445_403, w_445_404, 
  Loop Gates: I445_399.port1, I445_400.port1, I445_401.port2, I445_402.port2, I445_403.port1, 
  Loop Conditions: I445_399.port2=1, I445_400.port2=1, I445_401.port1=0, I445_402.port1=1, I445_403.port2=1, 
  (Singal Values: w_110_172=1, w_292_099=0, w_298_112=1, w_363_068=1, w_445_416=1, )

8)
  Loop Signals: w_445_402, w_445_408, w_445_409, w_445_410, w_445_411, w_445_412, w_445_413, w_445_414, w_445_416, 
  Loop Gates: I445_400.port2, I445_404.port2, I445_405.port1, I445_406.port1, I445_407.port2, I445_408.port2, I445_409.port2, I445_410.port1, I445_411.port2, 
  Loop Conditions: I445_400.port1=1, I445_404.port1=1, I445_405.port2=0, I445_407.port1=1, I445_408.port1=1, I445_409.port1=0, I445_411.port1=1, 
  (Singal Values: w_445_401=1, w_175_099=1, w_178_104=1, w_185_122=0, w_286_434=1, w_349_191=1, w_396_016=0, )

9)
  Loop Signals: w_186_061, w_186_062, w_186_063, w_186_064, w_186_065, w_186_066, w_186_067, w_186_068, 
  Loop Gates: I186_060.port1, I186_061.port1, I186_062.port1, I186_063.port1, I186_064.port2, I186_065.port2, I186_066.port1, I186_067.port1, 
  Loop Conditions: I186_060.port2=1, I186_061.port2=1, I186_063.port2=1, I186_064.port1=0, I186_065.port1=1, 
  (Singal Values: w_042_232=0, w_052_020=1, w_080_001=1, w_082_144=1, w_186_085=1, )

10)
  Loop Signals: w_186_065, w_186_072, w_186_073, w_186_074, w_186_075, w_186_076, w_186_077, w_186_078, w_186_079, w_186_080, w_186_081, w_186_082, w_186_083, w_186_085, 
  Loop Gates: I186_063.port2, I186_068.port1, I186_069.port2, I186_070.port2, I186_071.port2, I186_072.port1, I186_073.port1, I186_074.port2, I186_075.port1, I186_076.port2, I186_077.port1, I186_078.port2, I186_079.port1, I186_080.port2, 
  Loop Conditions: I186_063.port1=1, I186_068.port2=1, I186_069.port1=1, I186_070.port1=1, I186_071.port1=0, I186_072.port2=1, I186_073.port2=1, I186_074.port1=0, I186_075.port2=0, I186_076.port1=1, I186_077.port2=1, I186_078.port1=0, I186_080.port1=1, 
  (Singal Values: w_001_006=1, w_186_064=1, w_035_075=1, w_047_201=0, w_059_211=0, w_065_019=1, w_093_293=1, w_108_028=1, w_116_243=0, w_117_279=1, w_146_011=0, w_162_000=1, w_161_219=1, )

11)
  Loop Signals: w_088_456, w_088_460, w_088_461, w_088_462, w_088_463, w_088_464, w_088_465, w_088_466, w_088_467, w_088_468, w_088_469, w_088_471, 
  Loop Gates: I088_454.port2, I088_456.port2, I088_457.port2, I088_458.port2, I088_459.port1, I088_460.port2, I088_461.port1, I088_462.port1, I088_463.port1, I088_464.port2, I088_465.port1, I088_466.port2, 
  Loop Conditions: I088_454.port1=0, I088_456.port1=1, I088_457.port1=1, I088_458.port1=1, I088_459.port2=1, I088_460.port1=1, I088_461.port2=0, I088_462.port2=0, I088_463.port2=0, I088_464.port1=1, I088_466.port1=1, 
  (Singal Values: w_006_000=1, w_010_214=1, w_019_024=0, w_026_204=1, w_038_082=0, w_047_234=1, w_054_208=1, w_058_074=0, w_067_055=1, w_073_043=1, w_088_455=0, )

12)
  Loop Signals: w_372_147, w_372_148, w_372_149, w_372_150, w_372_151, w_372_152, w_372_153, w_372_154, 
  Loop Gates: I372_146.port1, I372_147.port1, I372_148.port1, I372_149.port2, I372_150.port2, I372_151.port1, I372_152.port1, I372_153.port1, 
  Loop Conditions: I372_146.port2=1, I372_147.port2=0, I372_148.port2=1, I372_149.port1=1, I372_150.port1=1, I372_151.port2=1, I372_152.port2=1, I372_153.port2=1, 
  (Singal Values: w_069_023=1, w_070_031=1, w_195_082=1, w_205_047=0, w_309_115=1, w_315_242=1, w_316_057=1, w_337_195=1, )

13)
  Loop Signals: w_484_092, w_484_093, w_484_094, w_484_095, w_484_096, 
  Loop Gates: I484_091.port1, I484_092.port1, I484_093.port1, I484_094.port1, I484_095.port1, 
  Loop Conditions: I484_091.port2=1, I484_092.port2=1, I484_094.port2=0, 
  (Singal Values: w_012_081=1, w_204_274=1, w_484_105=0, )

14)
  Loop Signals: w_203_367, w_203_368, w_203_369, w_203_370, w_203_371, w_203_372, w_203_373, 
  Loop Gates: I203_366.port1, I203_367.port2, I203_368.port1, I203_369.port1, I203_370.port2, I203_371.port1, I203_372.port1, 
  Loop Conditions: I203_367.port1=0, I203_368.port2=1, I203_369.port2=1, I203_370.port1=1, 
  (Singal Values: w_015_093=1, w_035_066=1, w_075_103=1, w_203_390=0, )

15)
  Loop Signals: w_138_241, w_138_242, w_138_243, w_138_244, w_138_245, w_138_246, w_138_247, w_138_248, 
  Loop Gates: I138_240.port1, I138_241.port2, I138_242.port2, I138_243.port1, I138_244.port1, I138_245.port1, I138_246.port1, I138_247.port1, 
  Loop Conditions: I138_240.port2=1, I138_241.port1=0, I138_242.port1=1, I138_243.port2=1, I138_244.port2=1, 
  (Singal Values: w_048_143=1, w_050_187=1, w_071_191=0, w_136_002=1, w_138_259=1, )

16)
  Loop Signals: w_138_244, w_138_252, w_138_253, w_138_254, w_138_255, w_138_256, w_138_257, w_138_259, 
  Loop Gates: I138_242.port1, I138_248.port1, I138_249.port2, I138_250.port2, I138_251.port1, I138_252.port1, I138_253.port1, I138_254.port2, 
  Loop Conditions: I138_242.port2=1, I138_248.port2=1, I138_249.port1=0, I138_250.port1=1, I138_251.port2=1, I138_252.port2=0, I138_254.port1=1, 
  (Singal Values: w_002_013=1, w_014_058=0, w_054_191=1, w_083_084=1, w_102_076=1, w_129_000=0, w_138_243=1, )

17)
  Loop Signals: w_039_500, w_039_513, w_039_514, w_039_515, w_039_516, w_039_517, w_039_518, w_039_519, w_039_520, w_039_522, 
  Loop Gates: I039_498.port2, I039_509.port1, I039_510.port2, I039_511.port1, I039_512.port1, I039_513.port1, I039_514.port2, I039_515.port1, I039_516.port1, I039_517.port2, 
  Loop Conditions: I039_498.port1=0, I039_510.port1=0, I039_512.port2=0, I039_513.port2=1, I039_514.port1=1, I039_517.port1=1, 
  (Singal Values: w_003_078=1, w_033_018=0, w_034_022=0, w_035_035=1, w_037_035=1, w_039_499=0, )

18)
  Loop Signals: w_226_396, w_226_397, w_226_398, w_226_399, w_226_400, w_226_401, w_226_402, w_226_403, 
  Loop Gates: I226_395.port1, I226_396.port1, I226_397.port2, I226_398.port1, I226_399.port1, I226_400.port1, I226_401.port1, I226_402.port1, 
  Loop Conditions: I226_395.port2=1, I226_397.port1=0, I226_400.port2=1, I226_401.port2=1, I226_402.port2=1, 
  (Singal Values: w_040_006=0, w_169_216=1, w_200_253=1, w_201_007=1, w_210_060=1, )

19)
  Loop Signals: w_317_341, w_317_342, w_317_343, w_317_344, w_317_345, w_317_346, w_317_347, w_317_348, w_317_349, w_317_350, w_317_351, 
  Loop Gates: I317_340.port2, I317_341.port1, I317_342.port1, I317_343.port1, I317_344.port2, I317_345.port2, I317_346.port1, I317_347.port1, I317_348.port2, I317_349.port1, I317_350.port1, 
  Loop Conditions: I317_340.port1=1, I317_342.port2=0, I317_343.port2=0, I317_344.port1=1, I317_345.port1=1, I317_346.port2=1, I317_348.port1=0, I317_349.port2=0, I317_350.port2=1, 
  (Singal Values: w_079_170=1, w_099_267=0, w_109_001=1, w_119_107=1, w_206_098=0, w_225_184=1, w_234_117=0, w_298_179=1, w_313_092=0, )

20)
  Loop Signals: w_303_197, w_303_198, w_303_199, w_303_200, 
  Loop Gates: I303_196.port2, I303_197.port1, I303_198.port2, I303_199.port1, 
  Loop Conditions: I303_196.port1=1, I303_198.port1=1, 
  (Singal Values: w_153_093=1, w_303_215=1, )

21)
  Loop Signals: w_303_198, w_303_204, w_303_205, w_303_206, w_303_207, w_303_208, w_303_209, w_303_210, w_303_211, w_303_212, w_303_213, w_303_215, 
  Loop Gates: I303_196.port1, I303_200.port1, I303_201.port1, I303_202.port1, I303_203.port1, I303_204.port1, I303_205.port1, I303_206.port1, I303_207.port2, I303_208.port1, I303_209.port1, I303_210.port2, 
  Loop Conditions: I303_196.port2=1, I303_202.port2=0, I303_203.port2=1, I303_205.port2=1, I303_207.port1=1, I303_208.port2=0, I303_210.port1=1, 
  (Singal Values: w_040_004=1, w_106_146=0, w_115_346=0, w_181_107=1, w_239_017=1, w_277_046=1, w_303_197=1, )

22)
  Loop Signals: w_318_385, w_318_394, w_318_395, w_318_396, w_318_397, w_318_398, w_318_399, w_318_401, 
  Loop Gates: I318_384.port2, I318_391.port2, I318_392.port1, I318_393.port1, I318_394.port2, I318_395.port1, I318_396.port1, I318_397.port2, 
  Loop Conditions: I318_384.port1=1, I318_391.port1=0, I318_393.port2=1, I318_394.port1=1, I318_395.port2=0, I318_397.port1=1, 
  (Singal Values: w_020_085=1, w_023_264=0, w_135_049=1, w_147_151=1, w_178_172=0, w_318_384=1, )

23)
  Loop Signals: w_375_267, w_375_276, w_375_277, w_375_278, w_375_279, w_375_280, w_375_281, w_375_282, w_375_283, w_375_284, w_375_285, w_375_286, w_375_288, 
  Loop Gates: I375_265.port1, I375_272.port2, I375_273.port1, I375_274.port2, I375_275.port1, I375_276.port2, I375_277.port2, I375_278.port1, I375_279.port1, I375_280.port2, I375_281.port2, I375_282.port1, I375_283.port2, 
  Loop Conditions: I375_265.port2=1, I375_272.port1=0, I375_274.port1=1, I375_276.port1=1, I375_277.port1=1, I375_278.port2=0, I375_279.port2=1, I375_280.port1=1, I375_281.port1=0, I375_283.port1=1, 
  (Singal Values: w_003_061=1, w_009_033=0, w_028_188=1, w_073_117=1, w_139_188=0, w_182_077=1, w_224_053=1, w_313_119=0, w_374_035=1, w_375_266=1, )

24)
  Loop Signals: w_093_429, w_093_434, w_093_435, w_093_436, w_093_437, w_093_438, w_093_439, w_093_440, w_093_441, w_093_442, w_093_443, w_093_444, w_093_445, w_093_447, 
  Loop Gates: I093_427.port1, I093_430.port1, I093_431.port1, I093_432.port1, I093_433.port1, I093_434.port2, I093_435.port2, I093_436.port1, I093_437.port1, I093_438.port2, I093_439.port2, I093_440.port1, I093_441.port1, I093_442.port2, 
  Loop Conditions: I093_427.port2=0, I093_430.port2=1, I093_432.port2=1, I093_433.port2=1, I093_434.port1=1, I093_435.port1=0, I093_436.port2=1, I093_438.port1=1, I093_439.port1=0, I093_442.port1=1, 
  (Singal Values: w_009_059=1, w_009_081=1, w_012_191=0, w_030_132=1, w_050_136=1, w_055_029=1, w_067_030=1, w_071_321=0, w_076_095=1, w_093_428=0, )

25)
  Loop Signals: w_127_507, w_127_508, w_127_509, w_127_510, w_127_511, w_127_512, w_127_513, w_127_514, w_127_515, w_127_516, w_127_517, 
  Loop Gates: I127_503.port2, I127_504.port2, I127_505.port1, I127_506.port2, I127_507.port2, I127_508.port2, I127_509.port1, I127_510.port2, I127_511.port2, I127_512.port1, I127_513.port1, 
  Loop Conditions: I127_503.port1=1, I127_504.port1=0, I127_506.port1=1, I127_507.port1=1, I127_508.port1=0, I127_510.port1=1, I127_511.port1=1, I127_512.port2=0, I127_513.port2=0, 
  (Singal Values: w_002_001=1, w_022_041=0, w_039_056=1, w_043_043=1, w_065_035=0, w_066_072=0, w_070_024=1, w_106_079=0, w_127_534=1, )

26)
  Loop Signals: w_022_164, w_022_165, w_022_166, w_022_167, w_022_168, w_022_169, w_022_170, w_022_171, w_022_172, w_022_173, 
  Loop Gates: I022_163.port2, I022_164.port1, I022_165.port1, I022_166.port1, I022_167.port2, I022_168.port2, I022_169.port1, I022_170.port2, I022_171.port2, I022_172.port2, 
  Loop Conditions: I022_163.port1=0, I022_164.port2=1, I022_165.port2=1, I022_166.port2=0, I022_167.port1=1, I022_168.port1=1, I022_169.port2=1, I022_170.port1=0, I022_171.port1=1, I022_172.port1=0, 
  (Singal Values: w_002_020=0, w_004_034=1, w_004_360=1, w_010_284=1, w_011_219=1, w_012_197=0, w_014_264=1, w_018_060=1, w_018_295=0, w_021_107=0, )

27)
  Loop Signals: w_173_283, w_173_284, w_173_285, w_173_286, w_173_287, w_173_288, w_173_289, w_173_290, w_173_291, w_173_292, 
  Loop Gates: I173_282.port1, I173_283.port1, I173_284.port2, I173_285.port2, I173_286.port1, I173_287.port2, I173_288.port1, I173_289.port2, I173_290.port1, I173_291.port2, 
  Loop Conditions: I173_284.port1=1, I173_285.port1=0, I173_286.port2=0, I173_287.port1=1, I173_288.port2=1, I173_289.port1=0, I173_290.port2=1, I173_291.port1=1, 
  (Singal Values: w_001_001=0, w_007_278=1, w_046_148=1, w_053_006=1, w_064_023=1, w_102_079=0, w_137_021=1, w_163_330=0, )

******* result_4.txt *********
1)
  Loop Breaker: w_139_230 

2)
  Loop Breaker: w_489_325 

3)
  Loop Breaker: w_158_039 

4)
  Loop Breaker: w_431_275 

5)
  Loop Breaker: w_029_256 

6)
  Loop Breaker: w_082_341 

7)
  Loop Breaker: w_445_402 

8)
  Loop Breaker: w_445_402 

9)
  Loop Breaker: w_186_065 

10)
  Loop Breaker: w_186_065 

11)
  Loop Breaker: w_088_456 

12)
  Loop Breaker: w_372_148 

13)
  Loop Breaker: w_484_096 

14)
  Loop Breaker: w_203_369 

15)
  Loop Breaker: w_138_244 

16)
  Loop Breaker: w_138_244 

17)
  Loop Breaker: w_039_500 

18)
  Loop Breaker: w_226_397 

19)
  Loop Breaker: w_317_342 

20)
  Loop Breaker: w_303_198 

21)
  Loop Breaker: w_303_198 

22)
  Loop Breaker: w_318_385 

23)
  Loop Breaker: w_375_267 

24)
  Loop Breaker: w_093_429 

25)
  Loop Breaker: w_127_515 

26)
  Loop Breaker: w_022_165 

27)
  Loop Breaker: w_173_284 

// ******* The results for this case End *********
*/
