// Gate Level Verilog Code Generated!
// GateLvl:40 GateNum:40 GateInputNum:2
// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_026, w_000_028, w_000_030, w_000_033, w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_026, w_000_028, w_000_030, w_000_033;
  output w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_026, w_000_028, w_000_030, w_000_033;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008;
  wire w_004_000, w_004_001, w_004_002, w_004_003, w_004_004, w_004_005, w_004_007, w_004_009, w_004_010;
  wire w_005_000, w_005_001, w_005_002, w_005_003, w_005_006, w_005_007, w_005_008, w_005_009, w_005_012, w_005_014, w_005_015, w_005_017, w_005_022, w_005_023, w_005_025, w_005_026;
  wire w_006_000, w_006_001, w_006_002;
  wire w_007_000, w_007_001, w_007_002, w_007_004, w_007_005, w_007_006, w_007_015, w_007_017, w_007_020, w_007_021, w_007_024, w_007_026, w_007_027, w_007_028, w_007_029, w_007_030, w_007_032, w_007_038, w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045;
  wire w_008_001, w_008_003, w_008_004, w_008_007, w_008_008, w_008_010, w_008_011, w_008_012;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_006, w_009_009, w_009_010;
  wire w_010_002, w_010_004, w_010_011, w_010_014, w_010_018, w_010_020, w_010_021, w_010_022, w_010_023, w_010_024, w_010_025, w_010_026, w_010_027;
  wire w_011_001, w_011_014, w_011_021, w_011_023, w_011_024, w_011_031, w_011_033;
  wire w_012_000, w_012_001, w_012_002, w_012_007, w_012_009;
  wire w_013_001, w_013_006;
  wire w_014_004, w_014_010, w_014_021;
  wire w_015_000;
  wire w_016_000, w_016_001, w_016_002;
  wire w_017_010;
  wire w_018_002, w_018_004, w_018_015, w_018_021;
  wire w_019_001;
  wire w_020_007, w_020_026, w_020_029, w_020_030, w_020_031, w_020_035, w_020_036, w_020_037, w_020_038, w_020_039, w_020_040, w_020_041, w_020_042, w_020_044;
  wire w_021_001, w_021_014, w_021_022, w_021_024;
  wire w_022_001, w_022_008, w_022_009;
  wire w_023_000, w_023_001;
  wire w_024_004;
  wire w_025_000;
  wire w_026_008;
  wire w_027_000;
  wire w_029_004, w_029_016, w_029_022;
  wire w_031_018, w_031_019, w_031_020, w_031_021, w_031_022, w_031_023, w_031_024, w_031_025, w_031_026, w_031_027, w_031_031, w_031_032, w_031_033, w_031_034, w_031_035, w_031_036, w_031_037, w_031_038, w_031_039, w_031_041;
  wire w_032_007;
  wire w_033_026, w_033_027, w_033_028, w_033_032, w_033_033, w_033_034, w_033_035, w_033_036, w_033_037, w_033_038, w_033_039, w_033_040;
  wire w_034_000;
  wire w_035_018, w_035_019, w_035_020, w_035_021, w_035_022, w_035_023, w_035_024, w_035_025, w_035_026, w_035_027, w_035_028;
  wire w_037_011;
  wire w_039_002;
  wire w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_002);
  nand2 I001_004(w_001_004, w_000_005, w_000_006);
  not1 I002_000(w_002_000, w_000_007);
  and2 I002_001(w_002_001, w_000_008, w_000_007);
  or2  I002_002(w_002_002, w_000_009, w_000_003);
  nand2 I002_003(w_002_003, w_001_004, w_000_010);
  not1 I002_004(w_002_004, w_001_002);
  or2  I002_005(w_002_005, w_000_011, w_000_012);
  or2  I002_006(w_002_006, w_001_004, w_000_013);
  not1 I002_007(w_002_007, w_000_014);
  or2  I003_000(w_003_000, w_001_001, w_002_004);
  or2  I003_001(w_003_001, w_002_002, w_001_001);
  or2  I003_002(w_003_002, w_000_004, w_000_015);
  or2  I003_003(w_003_003, w_001_004, w_001_002);
  and2 I003_004(w_003_004, w_000_016, w_000_014);
  nand2 I003_005(w_003_005, w_002_004, w_000_017);
  nand2 I003_006(w_003_006, w_000_018, w_002_004);
  and2 I003_007(w_003_007, w_000_011, w_002_007);
  and2 I003_008(w_003_008, w_000_019, w_001_001);
  not1 I004_000(w_004_000, w_003_008);
  not1 I004_001(w_004_001, w_002_002);
  nand2 I004_002(w_004_002, w_001_002, w_002_005);
  and2 I004_003(w_004_003, w_000_020, w_001_000);
  not1 I004_004(w_004_004, w_001_000);
  or2  I004_005(w_004_005, w_000_019, w_000_009);
  nand2 I004_007(w_004_007, w_001_002, w_003_007);
  and2 I004_009(w_004_009, w_000_021, w_000_022);
  nand2 I004_010(w_004_010, w_003_003, w_000_023);
  and2 I005_000(w_005_000, w_004_003, w_003_000);
  or2  I005_001(w_005_001, w_001_001, w_001_000);
  nand2 I005_002(w_005_002, w_003_004, w_003_001);
  not1 I005_003(w_005_003, w_003_002);
  nand2 I005_006(w_005_006, w_001_002, w_000_019);
  and2 I005_007(w_005_007, w_002_007, w_002_004);
  nand2 I005_008(w_005_008, w_002_002, w_001_003);
  nand2 I005_009(w_005_009, w_004_004, w_000_024);
  nand2 I005_012(w_005_012, w_003_004, w_003_006);
  or2  I005_014(w_005_014, w_002_005, w_001_004);
  nand2 I005_015(w_005_015, w_000_023, w_000_019);
  nand2 I005_017(w_005_017, w_004_004, w_004_002);
  nand2 I005_022(w_005_022, w_000_005, w_001_001);
  not1 I005_023(w_005_023, w_003_007);
  or2  I005_025(w_005_025, w_003_007, w_002_002);
  and2 I005_026(w_005_026, w_002_006, w_004_000);
  nand2 I006_000(w_006_000, w_003_002, w_003_001);
  or2  I006_001(w_006_001, w_002_004, w_003_003);
  or2  I006_002(w_006_002, w_005_008, w_003_004);
  and2 I007_000(w_007_000, w_005_015, w_004_004);
  and2 I007_001(w_007_001, w_003_001, w_004_005);
  not1 I007_002(w_007_002, w_004_005);
  and2 I007_004(w_007_004, w_001_002, w_000_009);
  and2 I007_005(w_007_005, w_002_006, w_001_001);
  or2  I007_006(w_007_006, w_006_000, w_004_004);
  not1 I007_015(w_007_015, w_002_004);
  nand2 I007_017(w_007_017, w_004_001, w_006_001);
  not1 I007_020(w_007_020, w_004_004);
  or2  I007_021(w_007_021, w_004_010, w_002_000);
  or2  I007_024(w_007_024, w_006_001, w_001_004);
  and2 I007_026(w_007_026, w_003_008, w_004_002);
  or2  I007_027(w_007_027, w_004_010, w_003_007);
  not1 I007_028(w_007_028, w_002_001);
  and2 I007_029(w_007_029, w_005_000, w_004_009);
  not1 I007_030(w_007_030, w_006_000);
  or2  I007_032(w_007_032, w_003_000, w_000_026);
  nand2 I007_038(w_007_038, w_002_001, w_002_002);
  or2  I007_039(w_007_041, w_007_040, w_006_000);
  nand2 I007_040(w_007_042, w_007_041, w_006_001);
  or2  I007_041(w_007_043, w_001_003, w_007_042);
  and2 I007_042(w_007_044, w_007_043, w_005_022);
  and2 I007_043(w_007_045, w_007_044, w_004_010);
  nand2 I007_044(w_007_040, w_001_001, w_007_045);
  nand2 I008_001(w_008_001, w_007_024, w_005_009);
  or2  I008_003(w_008_003, w_004_005, w_003_002);
  or2  I008_004(w_008_004, w_007_028, w_004_002);
  or2  I008_007(w_008_007, w_002_000, w_005_023);
  or2  I008_008(w_008_008, w_001_004, w_006_001);
  not1 I008_009(w_008_011, w_008_010);
  and2 I008_010(w_008_012, w_004_000, w_008_011);
  nand2 I008_011(w_008_010, w_006_000, w_008_012);
  nand2 I009_000(w_009_000, w_005_006, w_006_002);
  and2 I009_001(w_009_001, w_002_006, w_002_005);
  not1 I009_002(w_009_002, w_005_026);
  and2 I009_003(w_009_003, w_006_000, w_000_028);
  or2  I009_006(w_009_006, w_007_027, w_002_006);
  not1 I009_009(w_009_009, w_007_029);
  not1 I009_010(w_009_010, w_002_001);
  and2 I010_002(w_010_002, w_004_000, w_007_001);
  nand2 I010_004(w_010_004, w_009_003, w_002_002);
  nand2 I010_011(w_010_011, w_009_002, w_004_007);
  and2 I010_014(w_010_014, w_006_000, w_007_000);
  or2  I010_018(w_010_018, w_004_009, w_005_014);
  not1 I010_019(w_010_021, w_010_020);
  or2  I010_020(w_010_022, w_002_001, w_010_021);
  nand2 I010_021(w_010_023, w_010_022, w_001_000);
  and2 I010_022(w_010_024, w_007_032, w_010_023);
  and2 I010_023(w_010_025, w_009_001, w_010_024);
  and2 I010_024(w_010_026, w_010_025, w_007_002);
  not1 I010_025(w_010_027, w_010_026);
  not1 I010_026(w_010_020, w_010_027);
  or2  I011_001(w_011_001, w_002_005, w_003_004);
  nand2 I011_014(w_011_014, w_005_006, w_000_030);
  not1 I011_021(w_011_021, w_009_006);
  nand2 I011_023(w_011_023, w_006_001, w_005_002);
  nand2 I011_024(w_011_024, w_010_004, w_000_003);
  or2  I011_031(w_011_031, w_010_002, w_003_004);
  or2  I011_033(w_011_033, w_007_004, w_004_003);
  and2 I012_000(w_012_000, w_001_004, w_000_018);
  or2  I012_001(w_012_001, w_009_001, w_010_018);
  or2  I012_002(w_012_002, w_006_000, w_011_023);
  and2 I012_007(w_012_007, w_005_022, w_005_007);
  and2 I012_009(w_012_009, w_003_008, w_004_003);
  not1 I013_001(w_013_001, w_005_001);
  and2 I013_006(w_013_006, w_007_020, w_007_005);
  and2 I014_004(w_014_004, w_009_000, w_007_028);
  nand2 I014_010(w_014_010, w_003_003, w_010_018);
  or2  I014_021(w_014_021, w_011_001, w_008_003);
  not1 I015_000(w_015_000, w_005_025);
  or2  I016_000(w_016_000, w_015_000, w_014_021);
  nand2 I016_001(w_016_001, w_005_003, w_004_001);
  nand2 I016_002(w_016_002, w_011_024, w_000_033);
  or2  I017_010(w_017_010, w_011_014, w_004_002);
  and2 I018_002(w_018_002, w_001_002, w_004_001);
  and2 I018_004(w_018_004, w_015_000, w_000_019);
  nand2 I018_015(w_018_015, w_002_001, w_008_004);
  nand2 I018_021(w_018_021, w_001_003, w_002_003);
  and2 I019_001(w_019_001, w_007_006, w_015_000);
  not1 I020_007(w_020_007, w_009_003);
  nand2 I020_026(w_020_026, w_003_000, w_011_031);
  and2 I020_028(w_020_030, w_018_004, w_020_029);
  and2 I020_029(w_020_031, w_016_001, w_020_030);
  or2  I020_030(w_020_029, w_020_044, w_020_031);
  or2  I020_031(w_020_036, w_010_011, w_020_035);
  or2  I020_032(w_020_037, w_005_012, w_020_036);
  not1 I020_033(w_020_038, w_020_037);
  and2 I020_034(w_020_039, w_020_038, w_012_007);
  or2  I020_035(w_020_040, w_020_039, w_016_001);
  or2  I020_036(w_020_041, w_020_040, w_012_007);
  and2 I020_037(w_020_042, w_010_014, w_020_041);
  not1 I020_038(w_020_035, w_020_029);
  and2 I020_039(w_020_044, w_004_001, w_020_042);
  and2 I021_001(w_021_001, w_007_026, w_006_002);
  nand2 I021_014(w_021_014, w_000_008, w_014_010);
  or2  I021_022(w_021_022, w_012_009, w_014_004);
  or2  I021_024(w_021_024, w_019_001, w_016_000);
  nand2 I022_001(w_022_001, w_015_000, w_006_000);
  not1 I022_008(w_022_008, w_012_000);
  not1 I022_009(w_022_009, w_020_007);
  or2  I023_000(w_023_000, w_009_010, w_013_006);
  and2 I023_001(w_023_001, w_008_001, w_012_000);
  nand2 I024_004(w_024_004, w_023_000, w_022_008);
  or2  I025_000(w_025_000, w_007_015, w_002_004);
  not1 I026_008(w_026_008, w_012_002);
  not1 I027_000(w_027_000, w_007_017);
  not1 I029_004(w_029_004, w_003_004);
  and2 I029_016(w_029_016, w_011_033, w_021_022);
  or2  I029_022(w_029_022, w_022_001, w_024_004);
  nand2 I031_017(w_031_019, w_031_018, w_018_002);
  nand2 I031_018(w_031_020, w_031_019, w_004_003);
  or2  I031_019(w_031_021, w_031_020, w_013_001);
  not1 I031_020(w_031_022, w_031_021);
  not1 I031_021(w_031_023, w_031_022);
  not1 I031_022(w_031_024, w_031_023);
  nand2 I031_023(w_031_025, w_031_041, w_031_024);
  and2 I031_024(w_031_026, w_001_004, w_031_025);
  or2  I031_025(w_031_027, w_031_026, w_021_001);
  nand2 I031_026(w_031_018, w_031_027, w_004_010);
  nand2 I031_027(w_031_032, w_012_000, w_031_031);
  and2 I031_028(w_031_033, w_017_010, w_031_032);
  nand2 I031_029(w_031_034, w_031_033, w_027_000);
  and2 I031_030(w_031_035, w_025_000, w_031_034);
  and2 I031_031(w_031_036, w_005_000, w_031_035);
  not1 I031_032(w_031_037, w_031_036);
  and2 I031_033(w_031_038, w_023_001, w_031_037);
  and2 I031_034(w_031_039, w_008_008, w_031_038);
  not1 I031_035(w_031_031, w_031_025);
  and2 I031_036(w_031_041, w_027_000, w_031_039);
  or2  I032_007(w_032_007, w_002_001, w_023_001);
  and2 I033_025(w_033_027, w_033_026, w_008_007);
  and2 I033_026(w_033_028, w_007_030, w_033_027);
  and2 I033_027(w_033_026, w_016_000, w_033_028);
  and2 I033_028(w_033_033, w_033_032, w_023_001);
  and2 I033_029(w_033_034, w_033_033, w_029_016);
  or2  I033_030(w_033_035, w_033_034, w_001_000);
  not1 I033_031(w_033_036, w_033_035);
  not1 I033_032(w_033_037, w_033_036);
  and2 I033_033(w_033_038, w_033_037, w_011_021);
  or2  I033_034(w_033_039, w_014_021, w_033_038);
  and2 I033_035(w_033_040, w_033_039, w_021_014);
  not1 I033_036(w_033_032, w_033_040);
  and2 I034_000(w_034_000, w_018_021, w_007_038);
  and2 I035_017(w_035_019, w_005_026, w_035_018);
  and2 I035_018(w_035_020, w_035_019, w_008_007);
  not1 I035_019(w_035_021, w_035_020);
  nand2 I035_020(w_035_022, w_035_021, w_021_024);
  not1 I035_021(w_035_023, w_035_022);
  or2  I035_022(w_035_024, w_003_005, w_035_023);
  or2  I035_023(w_035_025, w_035_024, w_009_009);
  and2 I035_024(w_035_026, w_035_025, w_029_022);
  nand2 I035_025(w_035_027, w_026_008, w_035_026);
  and2 I035_026(w_035_028, w_005_017, w_035_027);
  nand2 I035_027(w_035_018, w_035_028, w_012_001);
  nand2 I037_011(w_037_011, w_023_001, w_020_026);
  and2 I039_002(w_039_002, w_006_000, w_034_000);
  or2  I040_000(w_040_000, w_004_005, w_018_015);
  or2  I040_001(w_040_001, w_029_004, w_016_002);
  or2  I040_002(w_040_002, w_000_015, w_039_002);
  and2 I040_003(w_040_003, w_006_000, w_001_003);
  nand2 I040_004(w_040_004, w_022_009, w_025_000);
  not1 I040_005(w_040_005, w_032_007);
  and2 I040_006(w_040_006, w_007_021, w_037_011);
  not1 I040_007(w_040_007, w_016_000);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_026, w_000_028, w_000_030, w_000_033, w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_026, w_000_028, w_000_030, w_000_033, w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
endmodule
*/
// ****** TestBench Module Defination End ******

/*
// ******* The results for this case *********
******* result_1.txt *********
1)
  Loop Signals: w_020_029, w_020_030, w_020_031, 
  Loop Gates: I020_028.port2, I020_029.port2, I020_030.port2, 

2)
  Loop Signals: w_020_029, w_020_035, w_020_036, w_020_037, w_020_038, w_020_039, w_020_040, w_020_041, w_020_042, w_020_044, 
  Loop Gates: I020_030.port1, I020_031.port2, I020_032.port2, I020_033.port1, I020_034.port1, I020_035.port1, I020_036.port1, I020_037.port2, I020_038.port1, I020_039.port2, 

3)
  Loop Signals: w_033_026, w_033_027, w_033_028, 
  Loop Gates: I033_025.port1, I033_026.port2, I033_027.port2, 

4)
  Loop Signals: w_035_018, w_035_019, w_035_020, w_035_021, w_035_022, w_035_023, w_035_024, w_035_025, w_035_026, w_035_027, w_035_028, 
  Loop Gates: I035_017.port2, I035_018.port1, I035_019.port1, I035_020.port1, I035_021.port1, I035_022.port2, I035_023.port1, I035_024.port1, I035_025.port2, I035_026.port2, I035_027.port1, 

5)
  Loop Signals: w_008_010, w_008_011, w_008_012, 
  Loop Gates: I008_009.port1, I008_010.port2, I008_011.port2, 

6)
  Loop Signals: w_031_018, w_031_019, w_031_020, w_031_021, w_031_022, w_031_023, w_031_024, w_031_025, w_031_026, w_031_027, 
  Loop Gates: I031_017.port1, I031_018.port1, I031_019.port1, I031_020.port1, I031_021.port1, I031_022.port1, I031_023.port2, I031_024.port2, I031_025.port1, I031_026.port1, 

7)
  Loop Signals: w_031_025, w_031_031, w_031_032, w_031_033, w_031_034, w_031_035, w_031_036, w_031_037, w_031_038, w_031_039, w_031_041, 
  Loop Gates: I031_023.port1, I031_027.port2, I031_028.port2, I031_029.port1, I031_030.port2, I031_031.port2, I031_032.port1, I031_033.port2, I031_034.port2, I031_035.port1, I031_036.port2, 

8)
  Loop Signals: w_010_020, w_010_021, w_010_022, w_010_023, w_010_024, w_010_025, w_010_026, w_010_027, 
  Loop Gates: I010_019.port1, I010_020.port2, I010_021.port1, I010_022.port2, I010_023.port2, I010_024.port1, I010_025.port1, I010_026.port1, 

9)
  Loop Signals: w_033_032, w_033_033, w_033_034, w_033_035, w_033_036, w_033_037, w_033_038, w_033_039, w_033_040, 
  Loop Gates: I033_028.port1, I033_029.port1, I033_030.port1, I033_031.port1, I033_032.port1, I033_033.port1, I033_034.port2, I033_035.port1, I033_036.port1, 

10)
  Loop Signals: w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045, 
  Loop Gates: I007_039.port1, I007_040.port1, I007_041.port2, I007_042.port1, I007_043.port1, I007_044.port2, 

******* result_2.txt *********
1)
  Loop Signals: w_020_029, w_020_030, w_020_031, 
  Loop Gates: I020_028.port2, I020_029.port2, I020_030.port2, 

2)
  Loop Signals: w_020_029, w_020_035, w_020_036, w_020_037, w_020_038, w_020_039, w_020_040, w_020_041, w_020_042, w_020_044, 
  Loop Gates: I020_030.port1, I020_031.port2, I020_032.port2, I020_033.port1, I020_034.port1, I020_035.port1, I020_036.port1, I020_037.port2, I020_038.port1, I020_039.port2, 

3)
  Loop Signals: w_033_026, w_033_027, w_033_028, 
  Loop Gates: I033_025.port1, I033_026.port2, I033_027.port2, 

4)
  Loop Signals: w_008_010, w_008_011, w_008_012, 
  Loop Gates: I008_009.port1, I008_010.port2, I008_011.port2, 

5)
  Loop Signals: w_010_020, w_010_021, w_010_022, w_010_023, w_010_024, w_010_025, w_010_026, w_010_027, 
  Loop Gates: I010_019.port1, I010_020.port2, I010_021.port1, I010_022.port2, I010_023.port2, I010_024.port1, I010_025.port1, I010_026.port1, 

6)
  Loop Signals: w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045, 
  Loop Gates: I007_039.port1, I007_040.port1, I007_041.port2, I007_042.port1, I007_043.port1, I007_044.port2, 

******* result_3.txt *********
1)
  Loop Signals: w_035_018, w_035_019, w_035_020, w_035_021, w_035_022, w_035_023, w_035_024, w_035_025, w_035_026, w_035_027, w_035_028, 
  Loop Gates: I035_017.port2, I035_018.port1, I035_019.port1, I035_020.port1, I035_021.port1, I035_022.port2, I035_023.port1, I035_024.port1, I035_025.port2, I035_026.port2, I035_027.port1, 
  Loop Conditions: I035_017.port1=1, I035_018.port2=1, I035_020.port2=1, I035_022.port1=0, I035_023.port2=0, I035_024.port2=1, I035_025.port1=1, I035_026.port1=1, I035_027.port2=1, 
  (Singal Values: w_003_005=0, w_005_017=1, w_005_026=1, w_008_007=1, w_009_009=0, w_012_001=1, w_021_024=1, w_026_008=1, w_029_022=1, )

2)
  Loop Signals: w_031_018, w_031_019, w_031_020, w_031_021, w_031_022, w_031_023, w_031_024, w_031_025, w_031_026, w_031_027, 
  Loop Gates: I031_017.port1, I031_018.port1, I031_019.port1, I031_020.port1, I031_021.port1, I031_022.port1, I031_023.port2, I031_024.port2, I031_025.port1, I031_026.port1, 
  Loop Conditions: I031_017.port2=1, I031_018.port2=1, I031_019.port2=0, I031_023.port1=1, I031_024.port1=1, I031_025.port2=0, I031_026.port2=1, 
  (Singal Values: w_001_004=1, w_004_003=1, w_004_010=1, w_013_001=0, w_018_002=1, w_021_001=0, w_031_041=1, )

3)
  Loop Signals: w_031_025, w_031_031, w_031_032, w_031_033, w_031_034, w_031_035, w_031_036, w_031_037, w_031_038, w_031_039, w_031_041, 
  Loop Gates: I031_023.port1, I031_027.port2, I031_028.port2, I031_029.port1, I031_030.port2, I031_031.port2, I031_032.port1, I031_033.port2, I031_034.port2, I031_035.port1, I031_036.port2, 
  Loop Conditions: I031_023.port2=1, I031_027.port1=1, I031_028.port1=1, I031_029.port2=1, I031_030.port1=1, I031_031.port1=1, I031_033.port1=1, I031_034.port1=1, I031_036.port1=1, 
  (Singal Values: w_005_000=1, w_008_008=1, w_012_000=1, w_017_010=1, w_023_001=1, w_025_000=1, w_027_000=1, w_031_024=1, )

4)
  Loop Signals: w_033_032, w_033_033, w_033_034, w_033_035, w_033_036, w_033_037, w_033_038, w_033_039, w_033_040, 
  Loop Gates: I033_028.port1, I033_029.port1, I033_030.port1, I033_031.port1, I033_032.port1, I033_033.port1, I033_034.port2, I033_035.port1, I033_036.port1, 
  Loop Conditions: I033_028.port2=1, I033_029.port2=1, I033_030.port2=0, I033_033.port2=1, I033_034.port1=0, I033_035.port2=1, 
  (Singal Values: w_001_000=0, w_011_021=1, w_014_021=0, w_021_014=1, w_023_001=1, w_029_016=1, )

******* result_4.txt *********
1)
  Loop Breaker: w_035_019 

2)
  Loop Breaker: w_031_025 

3)
  Loop Breaker: w_031_025 

4)
  Loop Breaker: w_033_033 

// ******* The results for this case End *********
*/
